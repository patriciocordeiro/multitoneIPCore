library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith;
use ieee.numeric_std.all;
use ieee.math_real.all;
entity moduloCounter is
	generic
	(
		--M:natural:= 2;
		fo: integer:= 1000000;
		fc: integer:= 100000000;
		N: integer:= 12; -- acumulator precision
		LTP:integer:= 8  --Look up table precision

	);
	port
	(
		clk: in std_logic;
		cnt: out std_logic_vector(N-1 downto 0);
		cntTrunc: out std_logic_vector(LTP-2 downto 0);
		MM: out unsigned(0 to N-1);
		mflag: out  std_logic;
		output : out  integer range -8192 to 8191;
		sinef : out  integer range -8192 to 8191;

		--sign_cnt: out integer range 0 to 2**N-1;
		firstIteration : out std_logic
	
	);
	end entity;
	architecture rtl of moduloCounter is
	
	constant temp:	integer range 0 to fc:= fc/fo;
	constant M: integer range 0 to (2**N)-1:= 2**N/temp+1;
	constant Mtrunc: integer range 0 to 300:=(M*(2**LTP))/2**N;
	--constant Mtrunc: integer range 0 to 300:=1;
	constant hN: unsigned(0 to N-1):= to_unsigned(2**(N-1), N);
	constant oneQtSize: unsigned (0 to LTP-1 ):= to_unsigned(2**(LTP-2),LTP); --one quater sine wave size
	constant acummToLutStep: integer range 0 to 2**(N-LTP):=2**(N-LTP); -- accumulator to lut step
	constant limit: unsigned(0 to N-1):=(to_unsigned(2**(N-1) ,N) + to_unsigned(2*acummToLutStep,N))/Mtrunc -1;
		
	
	signal cnt_temp: unsigned(0 to N-1):=to_unsigned(0,N);
	signal lutAddr: integer range 0 to 2**LTP-1;
	signal sine :integer range -8192 to 8191;
	signal sign_cnt_temp: integer range 0 to 2**N-1:=0;
	signal lutAddrM: integer range 0 to  2**LTP-1;
	signal fullLutAddr: integer range 0 to  2**N-1;
	--signal	sign_cnt: integer range 0 to 2**N-1:=0; 
	--signal c2tmp: unsigned (0 to LTP):=to_unsigned(0,N);

	
	begin
		process(clk, cnt_temp)
	 
	   variable flag: std_logic:='0';
	   variable firstIter: std_logic:='1'; -- signaling  the first iteration 
	   variable lutAddrPrev: integer range 0 to 2**LTP-1;
	  
		begin
		
		if rising_edge(clk) then
			----------------------------------------------------------------
			if (cnt_temp=0) then
			
				flag := '0'; --counter will increment 
					if (sign_cnt_temp < 2) then
					  sign_cnt_temp <= sign_cnt_temp + 1; --increment till first two positive sine quadrant
					else 
					  sign_cnt_temp <= 1;--restart the counter to one
					end if ;
			end if;
		 ----------------------------------------------------------------
		 ----$$$$$$$------------------------------------------------------------	
			if (cnt_temp>=0 AND (cnt_temp < limit) AND flag='0') then
			  --count while counter is greater than zero, limit not reached and counter increment
				--@@@@-------------------------------------------------
				if (firstIter = '0') then 
					--prevent the repetition of zero value
					cnt_temp<= cnt_temp + to_unsigned(acummToLutStep, N);
						--fullLutAddr<= to_integer(cnt_temp);
					firstIter :='1';
				else
					cnt_temp <= cnt_temp + 1;
					--fullLutAddr<= to_integer(cnt_temp);
				
					lutAddr <= to_integer(cnt_temp(0 to LTP-2));
				end if;
			   --@@@@--------------------------------------------------
			else
				flag:='1'; --  counter will decrement
					if (firstIter = '1') then 
					--prevent the repetition of zero value by jumping one step
						cnt_temp<= cnt_temp - to_unsigned(acummToLutStep, N);
						firstIter := '0'; 
							--fullLutAddr<= to_integer(cnt_temp);
					else
						cnt_temp <= cnt_temp - 1;
						lutAddr <= to_integer(cnt_temp(0 to LTP-2)); -- lookup table truncated counter
							--fullLutAddr<= to_integer(cnt_temp);
					end if;
			end if;
		----$$$$$$$------------------------------------------------------------	
				------------------------------
				if(lutAddrPrev/=lutAddr OR lutAddr=0) then
					lutAddrM <= lutAddr*Mtrunc;
					
				else
					lutAddrPrev := lutAddr;
				end if;
				------------------------------
				
				--&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
				--full counter
				if (fullLutAddr + M < (2**N-1)) then 
					fullLutAddr <= fullLutAddr + M;
				else 
					fullLutAddr <= 0;
				end if;
				--&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
				
		end if; --end rising_edge
		cnt <= std_logic_vector(cnt_temp);
		--cntTrunc <= std_logic_vector(cnt_temp(to_unsigned(N-LTP)));
		cntTrunc <= std_logic_vector(cnt_temp(0 to LTP-2));
		MM <= to_unsigned(M, N);
		mflag <= flag;
		--sign_cnt<= sign_cnt_temp;
		firstIteration <=firstIter;
  	end process;
  	
  	process(clk, lutAddrM)
		begin
	   if rising_edge(clk) then
			case lutAddrM is
 when 0 => sine <= 0;
 when 1 => sine <= 201;
 when 2 => sine <= 402;
 when 3 => sine <= 603;
 when 4 => sine <= 803;
 when 5 => sine <= 1003;
 when 6 => sine <= 1202;
 when 7 => sine <= 1400;
 when 8 => sine <= 1598;
 when 9 => sine <= 1795;
 when 10 => sine <= 1990;
 when 11 => sine <= 2185;
 when 12 => sine <= 2378;
 when 13 => sine <= 2569;
 when 14 => sine <= 2759;
 when 15 => sine <= 2948;
 when 16 => sine <= 3135;
 when 17 => sine <= 3319;
 when 18 => sine <= 3502;
 when 19 => sine <= 3683;
 when 20 => sine <= 3861;
 when 21 => sine <= 4037;
 when 22 => sine <= 4211;
 when 23 => sine <= 4382;
 when 24 => sine <= 4551;
 when 25 => sine <= 4716;
 when 26 => sine <= 4879;
 when 27 => sine <= 5039;
 when 28 => sine <= 5196;
 when 29 => sine <= 5350;
 when 30 => sine <= 5501;
 when 31 => sine <= 5648;
 when 32 => sine <= 5792;
 when 33 => sine <= 5932;
 when 34 => sine <= 6069;
 when 35 => sine <= 6202;
 when 36 => sine <= 6332;
 when 37 => sine <= 6457;
 when 38 => sine <= 6579;
 when 39 => sine <= 6697;
 when 40 => sine <= 6811;
 when 41 => sine <= 6920;
 when 42 => sine <= 7026;
 when 43 => sine <= 7127;
 when 44 => sine <= 7224;
 when 45 => sine <= 7316;
 when 46 => sine <= 7405;
 when 47 => sine <= 7488;
 when 48 => sine <= 7567;
 when 49 => sine <= 7642;
 when 50 => sine <= 7712;
 when 51 => sine <= 7778;
 when 52 => sine <= 7838;
 when 53 => sine <= 7894;
 when 54 => sine <= 7946;
 when 55 => sine <= 7992;
 when 56 => sine <= 8034;
 when 57 => sine <= 8070;
 when 58 => sine <= 8102;
 when 59 => sine <= 8129;
 when 60 => sine <= 8152;
 when 61 => sine <= 8169;
 when 62 => sine <= 8181;
 when 63 => sine <= 8189;
 when 64 => sine <= 8191;
 when 65 => sine <= 8189;
 when 66 => sine <= 8181;
 when 67 => sine <= 8169;
 when 68 => sine <= 8152;
 when 69 => sine <= 8129;
 when 70 => sine <= 8102;
 when 71 => sine <= 8070;
 when 72 => sine <= 8034;
 when 73 => sine <= 7992;
 when 74 => sine <= 7946;
 when 75 => sine <= 7894;
 when 76 => sine <= 7838;
 when 77 => sine <= 7778;
 when 78 => sine <= 7712;
 when 79 => sine <= 7642;
 when 80 => sine <= 7567;
 when 81 => sine <= 7488;
 when 82 => sine <= 7405;
 when 83 => sine <= 7316;
 when 84 => sine <= 7224;
 when 85 => sine <= 7127;
 when 86 => sine <= 7026;
 when 87 => sine <= 6920;
 when 88 => sine <= 6811;
 when 89 => sine <= 6697;
 when 90 => sine <= 6579;
 when 91 => sine <= 6457;
 when 92 => sine <= 6332;
 when 93 => sine <= 6202;
 when 94 => sine <= 6069;
 when 95 => sine <= 5932;
 when 96 => sine <= 5792;
 when 97 => sine <= 5648;
 when 98 => sine <= 5501;
 when 99 => sine <= 5350;
 when 100 => sine <= 5196;
 when 101 => sine <= 5039;
 when 102 => sine <= 4879;
 when 103 => sine <= 4716;
 when 104 => sine <= 4551;
 when 105 => sine <= 4382;
 when 106 => sine <= 4211;
 when 107 => sine <= 4037;
 when 108 => sine <= 3861;
 when 109 => sine <= 3683;
 when 110 => sine <= 3502;
 when 111 => sine <= 3319;
 when 112 => sine <= 3135;
 when 113 => sine <= 2948;
 when 114 => sine <= 2759;
 when 115 => sine <= 2569;
 when 116 => sine <= 2378;
 when 117 => sine <= 2185;
 when 118 => sine <= 1990;
 when 119 => sine <= 1795;
 when 120 => sine <= 1598;
 when 121 => sine <= 1400;
 when 122 => sine <= 1202;
 when 123 => sine <= 1003;
 when 124 => sine <= 803;
 when 125 => sine <= 603;
 when 126 => sine <= 402;
 when 127 => sine <= 201;
 when 128 => sine <= 0;
 when 129 => sine <= -201;
 when 130 => sine <= -402;
 when 131 => sine <= -603;
 when 132 => sine <= -803;
 when 133 => sine <= -1003;
 when 134 => sine <= -1202;
 when 135 => sine <= -1400;
 when 136 => sine <= -1598;
 when 137 => sine <= -1795;
 when 138 => sine <= -1990;
 when 139 => sine <= -2185;
 when 140 => sine <= -2378;
 when 141 => sine <= -2569;
 when 142 => sine <= -2759;
 when 143 => sine <= -2948;
 when 144 => sine <= -3135;
 when 145 => sine <= -3319;
 when 146 => sine <= -3502;
 when 147 => sine <= -3683;
 when 148 => sine <= -3861;
 when 149 => sine <= -4037;
 when 150 => sine <= -4211;
 when 151 => sine <= -4382;
 when 152 => sine <= -4551;
 when 153 => sine <= -4716;
 when 154 => sine <= -4879;
 when 155 => sine <= -5039;
 when 156 => sine <= -5196;
 when 157 => sine <= -5350;
 when 158 => sine <= -5501;
 when 159 => sine <= -5648;
 when 160 => sine <= -5792;
 when 161 => sine <= -5932;
 when 162 => sine <= -6069;
 when 163 => sine <= -6202;
 when 164 => sine <= -6332;
 when 165 => sine <= -6457;
 when 166 => sine <= -6579;
 when 167 => sine <= -6697;
 when 168 => sine <= -6811;
 when 169 => sine <= -6920;
 when 170 => sine <= -7026;
 when 171 => sine <= -7127;
 when 172 => sine <= -7224;
 when 173 => sine <= -7316;
 when 174 => sine <= -7405;
 when 175 => sine <= -7488;
 when 176 => sine <= -7567;
 when 177 => sine <= -7642;
 when 178 => sine <= -7712;
 when 179 => sine <= -7778;
 when 180 => sine <= -7838;
 when 181 => sine <= -7894;
 when 182 => sine <= -7946;
 when 183 => sine <= -7992;
 when 184 => sine <= -8034;
 when 185 => sine <= -8070;
 when 186 => sine <= -8102;
 when 187 => sine <= -8129;
 when 188 => sine <= -8152;
 when 189 => sine <= -8169;
 when 190 => sine <= -8181;
 when 191 => sine <= -8189;
 when 192 => sine <= -8191;
 when 193 => sine <= -8189;
 when 194 => sine <= -8181;
 when 195 => sine <= -8169;
 when 196 => sine <= -8152;
 when 197 => sine <= -8129;
 when 198 => sine <= -8102;
 when 199 => sine <= -8070;
 when 200 => sine <= -8034;
 when 201 => sine <= -7992;
 when 202 => sine <= -7946;
 when 203 => sine <= -7894;
 when 204 => sine <= -7838;
 when 205 => sine <= -7778;
 when 206 => sine <= -7712;
 when 207 => sine <= -7642;
 when 208 => sine <= -7567;
 when 209 => sine <= -7488;
 when 210 => sine <= -7405;
 when 211 => sine <= -7316;
 when 212 => sine <= -7224;
 when 213 => sine <= -7127;
 when 214 => sine <= -7026;
 when 215 => sine <= -6920;
 when 216 => sine <= -6811;
 when 217 => sine <= -6697;
 when 218 => sine <= -6579;
 when 219 => sine <= -6457;
 when 220 => sine <= -6332;
 when 221 => sine <= -6202;
 when 222 => sine <= -6069;
 when 223 => sine <= -5932;
 when 224 => sine <= -5792;
 when 225 => sine <= -5648;
 when 226 => sine <= -5501;
 when 227 => sine <= -5350;
 when 228 => sine <= -5196;
 when 229 => sine <= -5039;
 when 230 => sine <= -4879;
 when 231 => sine <= -4716;
 when 232 => sine <= -4551;
 when 233 => sine <= -4382;
 when 234 => sine <= -4211;
 when 235 => sine <= -4037;
 when 236 => sine <= -3861;
 when 237 => sine <= -3683;
 when 238 => sine <= -3502;
 when 239 => sine <= -3319;
 when 240 => sine <= -3135;
 when 241 => sine <= -2948;
 when 242 => sine <= -2759;
 when 243 => sine <= -2569;
 when 244 => sine <= -2378;
 when 245 => sine <= -2185;
 when 246 => sine <= -1990;
 when 247 => sine <= -1795;
 when 248 => sine <= -1598;
 when 249 => sine <= -1400;
 when 250 => sine <= -1202;
 when 251 => sine <= -1003;
 when 252 => sine <= -803;
 when 253 => sine <= -603;
 when 254 => sine <= -402;
 when 255 => sine <= -201;
 when others => sine <=0;
			end case;
		if (sign_cnt_temp < 2) then
        output <= sine;
    else
        output <= -sine;
    end if;
  
    end if;
	end process;

process(clk, fullLutAddr)
begin
	if rising_edge(clk) then
	 case fullLutAddr is
	 when 0 => sinef <= 0;
 when 1 => sinef <= 13;
 when 2 => sinef <= 25;
 when 3 => sinef <= 38;
 when 4 => sinef <= 50;
 when 5 => sinef <= 63;
 when 6 => sinef <= 75;
 when 7 => sinef <= 88;
 when 8 => sinef <= 101;
 when 9 => sinef <= 113;
 when 10 => sinef <= 126;
 when 11 => sinef <= 138;
 when 12 => sinef <= 151;
 when 13 => sinef <= 163;
 when 14 => sinef <= 176;
 when 15 => sinef <= 188;
 when 16 => sinef <= 201;
 when 17 => sinef <= 214;
 when 18 => sinef <= 226;
 when 19 => sinef <= 239;
 when 20 => sinef <= 251;
 when 21 => sinef <= 264;
 when 22 => sinef <= 276;
 when 23 => sinef <= 289;
 when 24 => sinef <= 301;
 when 25 => sinef <= 314;
 when 26 => sinef <= 327;
 when 27 => sinef <= 339;
 when 28 => sinef <= 352;
 when 29 => sinef <= 364;
 when 30 => sinef <= 377;
 when 31 => sinef <= 389;
 when 32 => sinef <= 402;
 when 33 => sinef <= 414;
 when 34 => sinef <= 427;
 when 35 => sinef <= 440;
 when 36 => sinef <= 452;
 when 37 => sinef <= 465;
 when 38 => sinef <= 477;
 when 39 => sinef <= 490;
 when 40 => sinef <= 502;
 when 41 => sinef <= 515;
 when 42 => sinef <= 527;
 when 43 => sinef <= 540;
 when 44 => sinef <= 552;
 when 45 => sinef <= 565;
 when 46 => sinef <= 578;
 when 47 => sinef <= 590;
 when 48 => sinef <= 603;
 when 49 => sinef <= 615;
 when 50 => sinef <= 628;
 when 51 => sinef <= 640;
 when 52 => sinef <= 653;
 when 53 => sinef <= 665;
 when 54 => sinef <= 678;
 when 55 => sinef <= 690;
 when 56 => sinef <= 703;
 when 57 => sinef <= 715;
 when 58 => sinef <= 728;
 when 59 => sinef <= 740;
 when 60 => sinef <= 753;
 when 61 => sinef <= 765;
 when 62 => sinef <= 778;
 when 63 => sinef <= 790;
 when 64 => sinef <= 803;
 when 65 => sinef <= 815;
 when 66 => sinef <= 828;
 when 67 => sinef <= 840;
 when 68 => sinef <= 853;
 when 69 => sinef <= 865;
 when 70 => sinef <= 878;
 when 71 => sinef <= 890;
 when 72 => sinef <= 903;
 when 73 => sinef <= 915;
 when 74 => sinef <= 928;
 when 75 => sinef <= 940;
 when 76 => sinef <= 953;
 when 77 => sinef <= 965;
 when 78 => sinef <= 978;
 when 79 => sinef <= 990;
 when 80 => sinef <= 1003;
 when 81 => sinef <= 1015;
 when 82 => sinef <= 1028;
 when 83 => sinef <= 1040;
 when 84 => sinef <= 1053;
 when 85 => sinef <= 1065;
 when 86 => sinef <= 1077;
 when 87 => sinef <= 1090;
 when 88 => sinef <= 1102;
 when 89 => sinef <= 1115;
 when 90 => sinef <= 1127;
 when 91 => sinef <= 1140;
 when 92 => sinef <= 1152;
 when 93 => sinef <= 1165;
 when 94 => sinef <= 1177;
 when 95 => sinef <= 1189;
 when 96 => sinef <= 1202;
 when 97 => sinef <= 1214;
 when 98 => sinef <= 1227;
 when 99 => sinef <= 1239;
 when 100 => sinef <= 1252;
 when 101 => sinef <= 1264;
 when 102 => sinef <= 1276;
 when 103 => sinef <= 1289;
 when 104 => sinef <= 1301;
 when 105 => sinef <= 1314;
 when 106 => sinef <= 1326;
 when 107 => sinef <= 1338;
 when 108 => sinef <= 1351;
 when 109 => sinef <= 1363;
 when 110 => sinef <= 1376;
 when 111 => sinef <= 1388;
 when 112 => sinef <= 1400;
 when 113 => sinef <= 1413;
 when 114 => sinef <= 1425;
 when 115 => sinef <= 1437;
 when 116 => sinef <= 1450;
 when 117 => sinef <= 1462;
 when 118 => sinef <= 1475;
 when 119 => sinef <= 1487;
 when 120 => sinef <= 1499;
 when 121 => sinef <= 1512;
 when 122 => sinef <= 1524;
 when 123 => sinef <= 1536;
 when 124 => sinef <= 1549;
 when 125 => sinef <= 1561;
 when 126 => sinef <= 1573;
 when 127 => sinef <= 1586;
 when 128 => sinef <= 1598;
 when 129 => sinef <= 1610;
 when 130 => sinef <= 1623;
 when 131 => sinef <= 1635;
 when 132 => sinef <= 1647;
 when 133 => sinef <= 1660;
 when 134 => sinef <= 1672;
 when 135 => sinef <= 1684;
 when 136 => sinef <= 1696;
 when 137 => sinef <= 1709;
 when 138 => sinef <= 1721;
 when 139 => sinef <= 1733;
 when 140 => sinef <= 1746;
 when 141 => sinef <= 1758;
 when 142 => sinef <= 1770;
 when 143 => sinef <= 1782;
 when 144 => sinef <= 1795;
 when 145 => sinef <= 1807;
 when 146 => sinef <= 1819;
 when 147 => sinef <= 1831;
 when 148 => sinef <= 1844;
 when 149 => sinef <= 1856;
 when 150 => sinef <= 1868;
 when 151 => sinef <= 1880;
 when 152 => sinef <= 1893;
 when 153 => sinef <= 1905;
 when 154 => sinef <= 1917;
 when 155 => sinef <= 1929;
 when 156 => sinef <= 1941;
 when 157 => sinef <= 1954;
 when 158 => sinef <= 1966;
 when 159 => sinef <= 1978;
 when 160 => sinef <= 1990;
 when 161 => sinef <= 2002;
 when 162 => sinef <= 2015;
 when 163 => sinef <= 2027;
 when 164 => sinef <= 2039;
 when 165 => sinef <= 2051;
 when 166 => sinef <= 2063;
 when 167 => sinef <= 2075;
 when 168 => sinef <= 2088;
 when 169 => sinef <= 2100;
 when 170 => sinef <= 2112;
 when 171 => sinef <= 2124;
 when 172 => sinef <= 2136;
 when 173 => sinef <= 2148;
 when 174 => sinef <= 2160;
 when 175 => sinef <= 2173;
 when 176 => sinef <= 2185;
 when 177 => sinef <= 2197;
 when 178 => sinef <= 2209;
 when 179 => sinef <= 2221;
 when 180 => sinef <= 2233;
 when 181 => sinef <= 2245;
 when 182 => sinef <= 2257;
 when 183 => sinef <= 2269;
 when 184 => sinef <= 2281;
 when 185 => sinef <= 2293;
 when 186 => sinef <= 2305;
 when 187 => sinef <= 2318;
 when 188 => sinef <= 2330;
 when 189 => sinef <= 2342;
 when 190 => sinef <= 2354;
 when 191 => sinef <= 2366;
 when 192 => sinef <= 2378;
 when 193 => sinef <= 2390;
 when 194 => sinef <= 2402;
 when 195 => sinef <= 2414;
 when 196 => sinef <= 2426;
 when 197 => sinef <= 2438;
 when 198 => sinef <= 2450;
 when 199 => sinef <= 2462;
 when 200 => sinef <= 2474;
 when 201 => sinef <= 2486;
 when 202 => sinef <= 2498;
 when 203 => sinef <= 2510;
 when 204 => sinef <= 2522;
 when 205 => sinef <= 2534;
 when 206 => sinef <= 2545;
 when 207 => sinef <= 2557;
 when 208 => sinef <= 2569;
 when 209 => sinef <= 2581;
 when 210 => sinef <= 2593;
 when 211 => sinef <= 2605;
 when 212 => sinef <= 2617;
 when 213 => sinef <= 2629;
 when 214 => sinef <= 2641;
 when 215 => sinef <= 2653;
 when 216 => sinef <= 2665;
 when 217 => sinef <= 2676;
 when 218 => sinef <= 2688;
 when 219 => sinef <= 2700;
 when 220 => sinef <= 2712;
 when 221 => sinef <= 2724;
 when 222 => sinef <= 2736;
 when 223 => sinef <= 2748;
 when 224 => sinef <= 2759;
 when 225 => sinef <= 2771;
 when 226 => sinef <= 2783;
 when 227 => sinef <= 2795;
 when 228 => sinef <= 2807;
 when 229 => sinef <= 2819;
 when 230 => sinef <= 2830;
 when 231 => sinef <= 2842;
 when 232 => sinef <= 2854;
 when 233 => sinef <= 2866;
 when 234 => sinef <= 2877;
 when 235 => sinef <= 2889;
 when 236 => sinef <= 2901;
 when 237 => sinef <= 2913;
 when 238 => sinef <= 2924;
 when 239 => sinef <= 2936;
 when 240 => sinef <= 2948;
 when 241 => sinef <= 2960;
 when 242 => sinef <= 2971;
 when 243 => sinef <= 2983;
 when 244 => sinef <= 2995;
 when 245 => sinef <= 3006;
 when 246 => sinef <= 3018;
 when 247 => sinef <= 3030;
 when 248 => sinef <= 3041;
 when 249 => sinef <= 3053;
 when 250 => sinef <= 3065;
 when 251 => sinef <= 3076;
 when 252 => sinef <= 3088;
 when 253 => sinef <= 3100;
 when 254 => sinef <= 3111;
 when 255 => sinef <= 3123;
 when 256 => sinef <= 3135;
 when 257 => sinef <= 3146;
 when 258 => sinef <= 3158;
 when 259 => sinef <= 3169;
 when 260 => sinef <= 3181;
 when 261 => sinef <= 3193;
 when 262 => sinef <= 3204;
 when 263 => sinef <= 3216;
 when 264 => sinef <= 3227;
 when 265 => sinef <= 3239;
 when 266 => sinef <= 3250;
 when 267 => sinef <= 3262;
 when 268 => sinef <= 3273;
 when 269 => sinef <= 3285;
 when 270 => sinef <= 3296;
 when 271 => sinef <= 3308;
 when 272 => sinef <= 3319;
 when 273 => sinef <= 3331;
 when 274 => sinef <= 3342;
 when 275 => sinef <= 3354;
 when 276 => sinef <= 3365;
 when 277 => sinef <= 3377;
 when 278 => sinef <= 3388;
 when 279 => sinef <= 3400;
 when 280 => sinef <= 3411;
 when 281 => sinef <= 3422;
 when 282 => sinef <= 3434;
 when 283 => sinef <= 3445;
 when 284 => sinef <= 3457;
 when 285 => sinef <= 3468;
 when 286 => sinef <= 3479;
 when 287 => sinef <= 3491;
 when 288 => sinef <= 3502;
 when 289 => sinef <= 3513;
 when 290 => sinef <= 3525;
 when 291 => sinef <= 3536;
 when 292 => sinef <= 3547;
 when 293 => sinef <= 3559;
 when 294 => sinef <= 3570;
 when 295 => sinef <= 3581;
 when 296 => sinef <= 3593;
 when 297 => sinef <= 3604;
 when 298 => sinef <= 3615;
 when 299 => sinef <= 3627;
 when 300 => sinef <= 3638;
 when 301 => sinef <= 3649;
 when 302 => sinef <= 3660;
 when 303 => sinef <= 3672;
 when 304 => sinef <= 3683;
 when 305 => sinef <= 3694;
 when 306 => sinef <= 3705;
 when 307 => sinef <= 3716;
 when 308 => sinef <= 3728;
 when 309 => sinef <= 3739;
 when 310 => sinef <= 3750;
 when 311 => sinef <= 3761;
 when 312 => sinef <= 3772;
 when 313 => sinef <= 3783;
 when 314 => sinef <= 3795;
 when 315 => sinef <= 3806;
 when 316 => sinef <= 3817;
 when 317 => sinef <= 3828;
 when 318 => sinef <= 3839;
 when 319 => sinef <= 3850;
 when 320 => sinef <= 3861;
 when 321 => sinef <= 3872;
 when 322 => sinef <= 3883;
 when 323 => sinef <= 3894;
 when 324 => sinef <= 3905;
 when 325 => sinef <= 3917;
 when 326 => sinef <= 3928;
 when 327 => sinef <= 3939;
 when 328 => sinef <= 3950;
 when 329 => sinef <= 3961;
 when 330 => sinef <= 3972;
 when 331 => sinef <= 3983;
 when 332 => sinef <= 3994;
 when 333 => sinef <= 4004;
 when 334 => sinef <= 4015;
 when 335 => sinef <= 4026;
 when 336 => sinef <= 4037;
 when 337 => sinef <= 4048;
 when 338 => sinef <= 4059;
 when 339 => sinef <= 4070;
 when 340 => sinef <= 4081;
 when 341 => sinef <= 4092;
 when 342 => sinef <= 4103;
 when 343 => sinef <= 4114;
 when 344 => sinef <= 4124;
 when 345 => sinef <= 4135;
 when 346 => sinef <= 4146;
 when 347 => sinef <= 4157;
 when 348 => sinef <= 4168;
 when 349 => sinef <= 4179;
 when 350 => sinef <= 4189;
 when 351 => sinef <= 4200;
 when 352 => sinef <= 4211;
 when 353 => sinef <= 4222;
 when 354 => sinef <= 4233;
 when 355 => sinef <= 4243;
 when 356 => sinef <= 4254;
 when 357 => sinef <= 4265;
 when 358 => sinef <= 4275;
 when 359 => sinef <= 4286;
 when 360 => sinef <= 4297;
 when 361 => sinef <= 4308;
 when 362 => sinef <= 4318;
 when 363 => sinef <= 4329;
 when 364 => sinef <= 4340;
 when 365 => sinef <= 4350;
 when 366 => sinef <= 4361;
 when 367 => sinef <= 4372;
 when 368 => sinef <= 4382;
 when 369 => sinef <= 4393;
 when 370 => sinef <= 4403;
 when 371 => sinef <= 4414;
 when 372 => sinef <= 4425;
 when 373 => sinef <= 4435;
 when 374 => sinef <= 4446;
 when 375 => sinef <= 4456;
 when 376 => sinef <= 4467;
 when 377 => sinef <= 4477;
 when 378 => sinef <= 4488;
 when 379 => sinef <= 4498;
 when 380 => sinef <= 4509;
 when 381 => sinef <= 4519;
 when 382 => sinef <= 4530;
 when 383 => sinef <= 4540;
 when 384 => sinef <= 4551;
 when 385 => sinef <= 4561;
 when 386 => sinef <= 4572;
 when 387 => sinef <= 4582;
 when 388 => sinef <= 4592;
 when 389 => sinef <= 4603;
 when 390 => sinef <= 4613;
 when 391 => sinef <= 4624;
 when 392 => sinef <= 4634;
 when 393 => sinef <= 4644;
 when 394 => sinef <= 4655;
 when 395 => sinef <= 4665;
 when 396 => sinef <= 4675;
 when 397 => sinef <= 4686;
 when 398 => sinef <= 4696;
 when 399 => sinef <= 4706;
 when 400 => sinef <= 4716;
 when 401 => sinef <= 4727;
 when 402 => sinef <= 4737;
 when 403 => sinef <= 4747;
 when 404 => sinef <= 4757;
 when 405 => sinef <= 4768;
 when 406 => sinef <= 4778;
 when 407 => sinef <= 4788;
 when 408 => sinef <= 4798;
 when 409 => sinef <= 4808;
 when 410 => sinef <= 4819;
 when 411 => sinef <= 4829;
 when 412 => sinef <= 4839;
 when 413 => sinef <= 4849;
 when 414 => sinef <= 4859;
 when 415 => sinef <= 4869;
 when 416 => sinef <= 4879;
 when 417 => sinef <= 4889;
 when 418 => sinef <= 4900;
 when 419 => sinef <= 4910;
 when 420 => sinef <= 4920;
 when 421 => sinef <= 4930;
 when 422 => sinef <= 4940;
 when 423 => sinef <= 4950;
 when 424 => sinef <= 4960;
 when 425 => sinef <= 4970;
 when 426 => sinef <= 4980;
 when 427 => sinef <= 4990;
 when 428 => sinef <= 5000;
 when 429 => sinef <= 5010;
 when 430 => sinef <= 5020;
 when 431 => sinef <= 5029;
 when 432 => sinef <= 5039;
 when 433 => sinef <= 5049;
 when 434 => sinef <= 5059;
 when 435 => sinef <= 5069;
 when 436 => sinef <= 5079;
 when 437 => sinef <= 5089;
 when 438 => sinef <= 5099;
 when 439 => sinef <= 5108;
 when 440 => sinef <= 5118;
 when 441 => sinef <= 5128;
 when 442 => sinef <= 5138;
 when 443 => sinef <= 5148;
 when 444 => sinef <= 5157;
 when 445 => sinef <= 5167;
 when 446 => sinef <= 5177;
 when 447 => sinef <= 5187;
 when 448 => sinef <= 5196;
 when 449 => sinef <= 5206;
 when 450 => sinef <= 5216;
 when 451 => sinef <= 5225;
 when 452 => sinef <= 5235;
 when 453 => sinef <= 5245;
 when 454 => sinef <= 5254;
 when 455 => sinef <= 5264;
 when 456 => sinef <= 5274;
 when 457 => sinef <= 5283;
 when 458 => sinef <= 5293;
 when 459 => sinef <= 5302;
 when 460 => sinef <= 5312;
 when 461 => sinef <= 5322;
 when 462 => sinef <= 5331;
 when 463 => sinef <= 5341;
 when 464 => sinef <= 5350;
 when 465 => sinef <= 5360;
 when 466 => sinef <= 5369;
 when 467 => sinef <= 5379;
 when 468 => sinef <= 5388;
 when 469 => sinef <= 5398;
 when 470 => sinef <= 5407;
 when 471 => sinef <= 5416;
 when 472 => sinef <= 5426;
 when 473 => sinef <= 5435;
 when 474 => sinef <= 5445;
 when 475 => sinef <= 5454;
 when 476 => sinef <= 5463;
 when 477 => sinef <= 5473;
 when 478 => sinef <= 5482;
 when 479 => sinef <= 5491;
 when 480 => sinef <= 5501;
 when 481 => sinef <= 5510;
 when 482 => sinef <= 5519;
 when 483 => sinef <= 5529;
 when 484 => sinef <= 5538;
 when 485 => sinef <= 5547;
 when 486 => sinef <= 5556;
 when 487 => sinef <= 5566;
 when 488 => sinef <= 5575;
 when 489 => sinef <= 5584;
 when 490 => sinef <= 5593;
 when 491 => sinef <= 5602;
 when 492 => sinef <= 5612;
 when 493 => sinef <= 5621;
 when 494 => sinef <= 5630;
 when 495 => sinef <= 5639;
 when 496 => sinef <= 5648;
 when 497 => sinef <= 5657;
 when 498 => sinef <= 5666;
 when 499 => sinef <= 5675;
 when 500 => sinef <= 5684;
 when 501 => sinef <= 5693;
 when 502 => sinef <= 5702;
 when 503 => sinef <= 5711;
 when 504 => sinef <= 5720;
 when 505 => sinef <= 5729;
 when 506 => sinef <= 5738;
 when 507 => sinef <= 5747;
 when 508 => sinef <= 5756;
 when 509 => sinef <= 5765;
 when 510 => sinef <= 5774;
 when 511 => sinef <= 5783;
 when 512 => sinef <= 5792;
 when 513 => sinef <= 5801;
 when 514 => sinef <= 5810;
 when 515 => sinef <= 5819;
 when 516 => sinef <= 5827;
 when 517 => sinef <= 5836;
 when 518 => sinef <= 5845;
 when 519 => sinef <= 5854;
 when 520 => sinef <= 5863;
 when 521 => sinef <= 5871;
 when 522 => sinef <= 5880;
 when 523 => sinef <= 5889;
 when 524 => sinef <= 5898;
 when 525 => sinef <= 5906;
 when 526 => sinef <= 5915;
 when 527 => sinef <= 5924;
 when 528 => sinef <= 5932;
 when 529 => sinef <= 5941;
 when 530 => sinef <= 5950;
 when 531 => sinef <= 5958;
 when 532 => sinef <= 5967;
 when 533 => sinef <= 5975;
 when 534 => sinef <= 5984;
 when 535 => sinef <= 5993;
 when 536 => sinef <= 6001;
 when 537 => sinef <= 6010;
 when 538 => sinef <= 6018;
 when 539 => sinef <= 6027;
 when 540 => sinef <= 6035;
 when 541 => sinef <= 6044;
 when 542 => sinef <= 6052;
 when 543 => sinef <= 6061;
 when 544 => sinef <= 6069;
 when 545 => sinef <= 6078;
 when 546 => sinef <= 6086;
 when 547 => sinef <= 6094;
 when 548 => sinef <= 6103;
 when 549 => sinef <= 6111;
 when 550 => sinef <= 6120;
 when 551 => sinef <= 6128;
 when 552 => sinef <= 6136;
 when 553 => sinef <= 6144;
 when 554 => sinef <= 6153;
 when 555 => sinef <= 6161;
 when 556 => sinef <= 6169;
 when 557 => sinef <= 6178;
 when 558 => sinef <= 6186;
 when 559 => sinef <= 6194;
 when 560 => sinef <= 6202;
 when 561 => sinef <= 6210;
 when 562 => sinef <= 6219;
 when 563 => sinef <= 6227;
 when 564 => sinef <= 6235;
 when 565 => sinef <= 6243;
 when 566 => sinef <= 6251;
 when 567 => sinef <= 6259;
 when 568 => sinef <= 6267;
 when 569 => sinef <= 6276;
 when 570 => sinef <= 6284;
 when 571 => sinef <= 6292;
 when 572 => sinef <= 6300;
 when 573 => sinef <= 6308;
 when 574 => sinef <= 6316;
 when 575 => sinef <= 6324;
 when 576 => sinef <= 6332;
 when 577 => sinef <= 6340;
 when 578 => sinef <= 6348;
 when 579 => sinef <= 6356;
 when 580 => sinef <= 6363;
 when 581 => sinef <= 6371;
 when 582 => sinef <= 6379;
 when 583 => sinef <= 6387;
 when 584 => sinef <= 6395;
 when 585 => sinef <= 6403;
 when 586 => sinef <= 6411;
 when 587 => sinef <= 6419;
 when 588 => sinef <= 6426;
 when 589 => sinef <= 6434;
 when 590 => sinef <= 6442;
 when 591 => sinef <= 6450;
 when 592 => sinef <= 6457;
 when 593 => sinef <= 6465;
 when 594 => sinef <= 6473;
 when 595 => sinef <= 6480;
 when 596 => sinef <= 6488;
 when 597 => sinef <= 6496;
 when 598 => sinef <= 6503;
 when 599 => sinef <= 6511;
 when 600 => sinef <= 6519;
 when 601 => sinef <= 6526;
 when 602 => sinef <= 6534;
 when 603 => sinef <= 6541;
 when 604 => sinef <= 6549;
 when 605 => sinef <= 6557;
 when 606 => sinef <= 6564;
 when 607 => sinef <= 6572;
 when 608 => sinef <= 6579;
 when 609 => sinef <= 6587;
 when 610 => sinef <= 6594;
 when 611 => sinef <= 6601;
 when 612 => sinef <= 6609;
 when 613 => sinef <= 6616;
 when 614 => sinef <= 6624;
 when 615 => sinef <= 6631;
 when 616 => sinef <= 6638;
 when 617 => sinef <= 6646;
 when 618 => sinef <= 6653;
 when 619 => sinef <= 6660;
 when 620 => sinef <= 6668;
 when 621 => sinef <= 6675;
 when 622 => sinef <= 6682;
 when 623 => sinef <= 6690;
 when 624 => sinef <= 6697;
 when 625 => sinef <= 6704;
 when 626 => sinef <= 6711;
 when 627 => sinef <= 6718;
 when 628 => sinef <= 6726;
 when 629 => sinef <= 6733;
 when 630 => sinef <= 6740;
 when 631 => sinef <= 6747;
 when 632 => sinef <= 6754;
 when 633 => sinef <= 6761;
 when 634 => sinef <= 6768;
 when 635 => sinef <= 6775;
 when 636 => sinef <= 6783;
 when 637 => sinef <= 6790;
 when 638 => sinef <= 6797;
 when 639 => sinef <= 6804;
 when 640 => sinef <= 6811;
 when 641 => sinef <= 6818;
 when 642 => sinef <= 6824;
 when 643 => sinef <= 6831;
 when 644 => sinef <= 6838;
 when 645 => sinef <= 6845;
 when 646 => sinef <= 6852;
 when 647 => sinef <= 6859;
 when 648 => sinef <= 6866;
 when 649 => sinef <= 6873;
 when 650 => sinef <= 6880;
 when 651 => sinef <= 6886;
 when 652 => sinef <= 6893;
 when 653 => sinef <= 6900;
 when 654 => sinef <= 6907;
 when 655 => sinef <= 6913;
 when 656 => sinef <= 6920;
 when 657 => sinef <= 6927;
 when 658 => sinef <= 6934;
 when 659 => sinef <= 6940;
 when 660 => sinef <= 6947;
 when 661 => sinef <= 6954;
 when 662 => sinef <= 6960;
 when 663 => sinef <= 6967;
 when 664 => sinef <= 6973;
 when 665 => sinef <= 6980;
 when 666 => sinef <= 6987;
 when 667 => sinef <= 6993;
 when 668 => sinef <= 7000;
 when 669 => sinef <= 7006;
 when 670 => sinef <= 7013;
 when 671 => sinef <= 7019;
 when 672 => sinef <= 7026;
 when 673 => sinef <= 7032;
 when 674 => sinef <= 7039;
 when 675 => sinef <= 7045;
 when 676 => sinef <= 7051;
 when 677 => sinef <= 7058;
 when 678 => sinef <= 7064;
 when 679 => sinef <= 7070;
 when 680 => sinef <= 7077;
 when 681 => sinef <= 7083;
 when 682 => sinef <= 7089;
 when 683 => sinef <= 7096;
 when 684 => sinef <= 7102;
 when 685 => sinef <= 7108;
 when 686 => sinef <= 7114;
 when 687 => sinef <= 7121;
 when 688 => sinef <= 7127;
 when 689 => sinef <= 7133;
 when 690 => sinef <= 7139;
 when 691 => sinef <= 7145;
 when 692 => sinef <= 7152;
 when 693 => sinef <= 7158;
 when 694 => sinef <= 7164;
 when 695 => sinef <= 7170;
 when 696 => sinef <= 7176;
 when 697 => sinef <= 7182;
 when 698 => sinef <= 7188;
 when 699 => sinef <= 7194;
 when 700 => sinef <= 7200;
 when 701 => sinef <= 7206;
 when 702 => sinef <= 7212;
 when 703 => sinef <= 7218;
 when 704 => sinef <= 7224;
 when 705 => sinef <= 7230;
 when 706 => sinef <= 7236;
 when 707 => sinef <= 7242;
 when 708 => sinef <= 7247;
 when 709 => sinef <= 7253;
 when 710 => sinef <= 7259;
 when 711 => sinef <= 7265;
 when 712 => sinef <= 7271;
 when 713 => sinef <= 7276;
 when 714 => sinef <= 7282;
 when 715 => sinef <= 7288;
 when 716 => sinef <= 7294;
 when 717 => sinef <= 7299;
 when 718 => sinef <= 7305;
 when 719 => sinef <= 7311;
 when 720 => sinef <= 7316;
 when 721 => sinef <= 7322;
 when 722 => sinef <= 7328;
 when 723 => sinef <= 7333;
 when 724 => sinef <= 7339;
 when 725 => sinef <= 7344;
 when 726 => sinef <= 7350;
 when 727 => sinef <= 7356;
 when 728 => sinef <= 7361;
 when 729 => sinef <= 7367;
 when 730 => sinef <= 7372;
 when 731 => sinef <= 7377;
 when 732 => sinef <= 7383;
 when 733 => sinef <= 7388;
 when 734 => sinef <= 7394;
 when 735 => sinef <= 7399;
 when 736 => sinef <= 7405;
 when 737 => sinef <= 7410;
 when 738 => sinef <= 7415;
 when 739 => sinef <= 7421;
 when 740 => sinef <= 7426;
 when 741 => sinef <= 7431;
 when 742 => sinef <= 7436;
 when 743 => sinef <= 7442;
 when 744 => sinef <= 7447;
 when 745 => sinef <= 7452;
 when 746 => sinef <= 7457;
 when 747 => sinef <= 7463;
 when 748 => sinef <= 7468;
 when 749 => sinef <= 7473;
 when 750 => sinef <= 7478;
 when 751 => sinef <= 7483;
 when 752 => sinef <= 7488;
 when 753 => sinef <= 7493;
 when 754 => sinef <= 7498;
 when 755 => sinef <= 7503;
 when 756 => sinef <= 7509;
 when 757 => sinef <= 7514;
 when 758 => sinef <= 7519;
 when 759 => sinef <= 7524;
 when 760 => sinef <= 7528;
 when 761 => sinef <= 7533;
 when 762 => sinef <= 7538;
 when 763 => sinef <= 7543;
 when 764 => sinef <= 7548;
 when 765 => sinef <= 7553;
 when 766 => sinef <= 7558;
 when 767 => sinef <= 7563;
 when 768 => sinef <= 7567;
 when 769 => sinef <= 7572;
 when 770 => sinef <= 7577;
 when 771 => sinef <= 7582;
 when 772 => sinef <= 7587;
 when 773 => sinef <= 7591;
 when 774 => sinef <= 7596;
 when 775 => sinef <= 7601;
 when 776 => sinef <= 7605;
 when 777 => sinef <= 7610;
 when 778 => sinef <= 7615;
 when 779 => sinef <= 7619;
 when 780 => sinef <= 7624;
 when 781 => sinef <= 7628;
 when 782 => sinef <= 7633;
 when 783 => sinef <= 7638;
 when 784 => sinef <= 7642;
 when 785 => sinef <= 7647;
 when 786 => sinef <= 7651;
 when 787 => sinef <= 7656;
 when 788 => sinef <= 7660;
 when 789 => sinef <= 7665;
 when 790 => sinef <= 7669;
 when 791 => sinef <= 7673;
 when 792 => sinef <= 7678;
 when 793 => sinef <= 7682;
 when 794 => sinef <= 7686;
 when 795 => sinef <= 7691;
 when 796 => sinef <= 7695;
 when 797 => sinef <= 7699;
 when 798 => sinef <= 7704;
 when 799 => sinef <= 7708;
 when 800 => sinef <= 7712;
 when 801 => sinef <= 7716;
 when 802 => sinef <= 7721;
 when 803 => sinef <= 7725;
 when 804 => sinef <= 7729;
 when 805 => sinef <= 7733;
 when 806 => sinef <= 7737;
 when 807 => sinef <= 7741;
 when 808 => sinef <= 7745;
 when 809 => sinef <= 7750;
 when 810 => sinef <= 7754;
 when 811 => sinef <= 7758;
 when 812 => sinef <= 7762;
 when 813 => sinef <= 7766;
 when 814 => sinef <= 7770;
 when 815 => sinef <= 7774;
 when 816 => sinef <= 7778;
 when 817 => sinef <= 7782;
 when 818 => sinef <= 7785;
 when 819 => sinef <= 7789;
 when 820 => sinef <= 7793;
 when 821 => sinef <= 7797;
 when 822 => sinef <= 7801;
 when 823 => sinef <= 7805;
 when 824 => sinef <= 7809;
 when 825 => sinef <= 7812;
 when 826 => sinef <= 7816;
 when 827 => sinef <= 7820;
 when 828 => sinef <= 7824;
 when 829 => sinef <= 7827;
 when 830 => sinef <= 7831;
 when 831 => sinef <= 7835;
 when 832 => sinef <= 7838;
 when 833 => sinef <= 7842;
 when 834 => sinef <= 7846;
 when 835 => sinef <= 7849;
 when 836 => sinef <= 7853;
 when 837 => sinef <= 7856;
 when 838 => sinef <= 7860;
 when 839 => sinef <= 7863;
 when 840 => sinef <= 7867;
 when 841 => sinef <= 7870;
 when 842 => sinef <= 7874;
 when 843 => sinef <= 7877;
 when 844 => sinef <= 7881;
 when 845 => sinef <= 7884;
 when 846 => sinef <= 7888;
 when 847 => sinef <= 7891;
 when 848 => sinef <= 7894;
 when 849 => sinef <= 7898;
 when 850 => sinef <= 7901;
 when 851 => sinef <= 7904;
 when 852 => sinef <= 7908;
 when 853 => sinef <= 7911;
 when 854 => sinef <= 7914;
 when 855 => sinef <= 7917;
 when 856 => sinef <= 7921;
 when 857 => sinef <= 7924;
 when 858 => sinef <= 7927;
 when 859 => sinef <= 7930;
 when 860 => sinef <= 7933;
 when 861 => sinef <= 7936;
 when 862 => sinef <= 7939;
 when 863 => sinef <= 7942;
 when 864 => sinef <= 7946;
 when 865 => sinef <= 7949;
 when 866 => sinef <= 7952;
 when 867 => sinef <= 7955;
 when 868 => sinef <= 7958;
 when 869 => sinef <= 7961;
 when 870 => sinef <= 7964;
 when 871 => sinef <= 7966;
 when 872 => sinef <= 7969;
 when 873 => sinef <= 7972;
 when 874 => sinef <= 7975;
 when 875 => sinef <= 7978;
 when 876 => sinef <= 7981;
 when 877 => sinef <= 7984;
 when 878 => sinef <= 7986;
 when 879 => sinef <= 7989;
 when 880 => sinef <= 7992;
 when 881 => sinef <= 7995;
 when 882 => sinef <= 7997;
 when 883 => sinef <= 8000;
 when 884 => sinef <= 8003;
 when 885 => sinef <= 8006;
 when 886 => sinef <= 8008;
 when 887 => sinef <= 8011;
 when 888 => sinef <= 8013;
 when 889 => sinef <= 8016;
 when 890 => sinef <= 8019;
 when 891 => sinef <= 8021;
 when 892 => sinef <= 8024;
 when 893 => sinef <= 8026;
 when 894 => sinef <= 8029;
 when 895 => sinef <= 8031;
 when 896 => sinef <= 8034;
 when 897 => sinef <= 8036;
 when 898 => sinef <= 8038;
 when 899 => sinef <= 8041;
 when 900 => sinef <= 8043;
 when 901 => sinef <= 8046;
 when 902 => sinef <= 8048;
 when 903 => sinef <= 8050;
 when 904 => sinef <= 8053;
 when 905 => sinef <= 8055;
 when 906 => sinef <= 8057;
 when 907 => sinef <= 8059;
 when 908 => sinef <= 8062;
 when 909 => sinef <= 8064;
 when 910 => sinef <= 8066;
 when 911 => sinef <= 8068;
 when 912 => sinef <= 8070;
 when 913 => sinef <= 8073;
 when 914 => sinef <= 8075;
 when 915 => sinef <= 8077;
 when 916 => sinef <= 8079;
 when 917 => sinef <= 8081;
 when 918 => sinef <= 8083;
 when 919 => sinef <= 8085;
 when 920 => sinef <= 8087;
 when 921 => sinef <= 8089;
 when 922 => sinef <= 8091;
 when 923 => sinef <= 8093;
 when 924 => sinef <= 8095;
 when 925 => sinef <= 8097;
 when 926 => sinef <= 8099;
 when 927 => sinef <= 8100;
 when 928 => sinef <= 8102;
 when 929 => sinef <= 8104;
 when 930 => sinef <= 8106;
 when 931 => sinef <= 8108;
 when 932 => sinef <= 8110;
 when 933 => sinef <= 8111;
 when 934 => sinef <= 8113;
 when 935 => sinef <= 8115;
 when 936 => sinef <= 8116;
 when 937 => sinef <= 8118;
 when 938 => sinef <= 8120;
 when 939 => sinef <= 8121;
 when 940 => sinef <= 8123;
 when 941 => sinef <= 8125;
 when 942 => sinef <= 8126;
 when 943 => sinef <= 8128;
 when 944 => sinef <= 8129;
 when 945 => sinef <= 8131;
 when 946 => sinef <= 8132;
 when 947 => sinef <= 8134;
 when 948 => sinef <= 8135;
 when 949 => sinef <= 8137;
 when 950 => sinef <= 8138;
 when 951 => sinef <= 8140;
 when 952 => sinef <= 8141;
 when 953 => sinef <= 8142;
 when 954 => sinef <= 8144;
 when 955 => sinef <= 8145;
 when 956 => sinef <= 8146;
 when 957 => sinef <= 8148;
 when 958 => sinef <= 8149;
 when 959 => sinef <= 8150;
 when 960 => sinef <= 8152;
 when 961 => sinef <= 8153;
 when 962 => sinef <= 8154;
 when 963 => sinef <= 8155;
 when 964 => sinef <= 8156;
 when 965 => sinef <= 8157;
 when 966 => sinef <= 8159;
 when 967 => sinef <= 8160;
 when 968 => sinef <= 8161;
 when 969 => sinef <= 8162;
 when 970 => sinef <= 8163;
 when 971 => sinef <= 8164;
 when 972 => sinef <= 8165;
 when 973 => sinef <= 8166;
 when 974 => sinef <= 8167;
 when 975 => sinef <= 8168;
 when 976 => sinef <= 8169;
 when 977 => sinef <= 8170;
 when 978 => sinef <= 8171;
 when 979 => sinef <= 8171;
 when 980 => sinef <= 8172;
 when 981 => sinef <= 8173;
 when 982 => sinef <= 8174;
 when 983 => sinef <= 8175;
 when 984 => sinef <= 8176;
 when 985 => sinef <= 8176;
 when 986 => sinef <= 8177;
 when 987 => sinef <= 8178;
 when 988 => sinef <= 8179;
 when 989 => sinef <= 8179;
 when 990 => sinef <= 8180;
 when 991 => sinef <= 8181;
 when 992 => sinef <= 8181;
 when 993 => sinef <= 8182;
 when 994 => sinef <= 8182;
 when 995 => sinef <= 8183;
 when 996 => sinef <= 8183;
 when 997 => sinef <= 8184;
 when 998 => sinef <= 8184;
 when 999 => sinef <= 8185;
 when 1000 => sinef <= 8185;
 when 1001 => sinef <= 8186;
 when 1002 => sinef <= 8186;
 when 1003 => sinef <= 8187;
 when 1004 => sinef <= 8187;
 when 1005 => sinef <= 8188;
 when 1006 => sinef <= 8188;
 when 1007 => sinef <= 8188;
 when 1008 => sinef <= 8189;
 when 1009 => sinef <= 8189;
 when 1010 => sinef <= 8189;
 when 1011 => sinef <= 8189;
 when 1012 => sinef <= 8190;
 when 1013 => sinef <= 8190;
 when 1014 => sinef <= 8190;
 when 1015 => sinef <= 8190;
 when 1016 => sinef <= 8190;
 when 1017 => sinef <= 8191;
 when 1018 => sinef <= 8191;
 when 1019 => sinef <= 8191;
 when 1020 => sinef <= 8191;
 when 1021 => sinef <= 8191;
 when 1022 => sinef <= 8191;
 when 1023 => sinef <= 8191;
 when 1024 => sinef <= 8191;
 when 1025 => sinef <= 8191;
 when 1026 => sinef <= 8191;
 when 1027 => sinef <= 8191;
 when 1028 => sinef <= 8191;
 when 1029 => sinef <= 8191;
 when 1030 => sinef <= 8191;
 when 1031 => sinef <= 8191;
 when 1032 => sinef <= 8190;
 when 1033 => sinef <= 8190;
 when 1034 => sinef <= 8190;
 when 1035 => sinef <= 8190;
 when 1036 => sinef <= 8190;
 when 1037 => sinef <= 8189;
 when 1038 => sinef <= 8189;
 when 1039 => sinef <= 8189;
 when 1040 => sinef <= 8189;
 when 1041 => sinef <= 8188;
 when 1042 => sinef <= 8188;
 when 1043 => sinef <= 8188;
 when 1044 => sinef <= 8187;
 when 1045 => sinef <= 8187;
 when 1046 => sinef <= 8186;
 when 1047 => sinef <= 8186;
 when 1048 => sinef <= 8185;
 when 1049 => sinef <= 8185;
 when 1050 => sinef <= 8184;
 when 1051 => sinef <= 8184;
 when 1052 => sinef <= 8183;
 when 1053 => sinef <= 8183;
 when 1054 => sinef <= 8182;
 when 1055 => sinef <= 8182;
 when 1056 => sinef <= 8181;
 when 1057 => sinef <= 8181;
 when 1058 => sinef <= 8180;
 when 1059 => sinef <= 8179;
 when 1060 => sinef <= 8179;
 when 1061 => sinef <= 8178;
 when 1062 => sinef <= 8177;
 when 1063 => sinef <= 8176;
 when 1064 => sinef <= 8176;
 when 1065 => sinef <= 8175;
 when 1066 => sinef <= 8174;
 when 1067 => sinef <= 8173;
 when 1068 => sinef <= 8172;
 when 1069 => sinef <= 8171;
 when 1070 => sinef <= 8171;
 when 1071 => sinef <= 8170;
 when 1072 => sinef <= 8169;
 when 1073 => sinef <= 8168;
 when 1074 => sinef <= 8167;
 when 1075 => sinef <= 8166;
 when 1076 => sinef <= 8165;
 when 1077 => sinef <= 8164;
 when 1078 => sinef <= 8163;
 when 1079 => sinef <= 8162;
 when 1080 => sinef <= 8161;
 when 1081 => sinef <= 8160;
 when 1082 => sinef <= 8159;
 when 1083 => sinef <= 8157;
 when 1084 => sinef <= 8156;
 when 1085 => sinef <= 8155;
 when 1086 => sinef <= 8154;
 when 1087 => sinef <= 8153;
 when 1088 => sinef <= 8152;
 when 1089 => sinef <= 8150;
 when 1090 => sinef <= 8149;
 when 1091 => sinef <= 8148;
 when 1092 => sinef <= 8146;
 when 1093 => sinef <= 8145;
 when 1094 => sinef <= 8144;
 when 1095 => sinef <= 8142;
 when 1096 => sinef <= 8141;
 when 1097 => sinef <= 8140;
 when 1098 => sinef <= 8138;
 when 1099 => sinef <= 8137;
 when 1100 => sinef <= 8135;
 when 1101 => sinef <= 8134;
 when 1102 => sinef <= 8132;
 when 1103 => sinef <= 8131;
 when 1104 => sinef <= 8129;
 when 1105 => sinef <= 8128;
 when 1106 => sinef <= 8126;
 when 1107 => sinef <= 8125;
 when 1108 => sinef <= 8123;
 when 1109 => sinef <= 8121;
 when 1110 => sinef <= 8120;
 when 1111 => sinef <= 8118;
 when 1112 => sinef <= 8116;
 when 1113 => sinef <= 8115;
 when 1114 => sinef <= 8113;
 when 1115 => sinef <= 8111;
 when 1116 => sinef <= 8110;
 when 1117 => sinef <= 8108;
 when 1118 => sinef <= 8106;
 when 1119 => sinef <= 8104;
 when 1120 => sinef <= 8102;
 when 1121 => sinef <= 8100;
 when 1122 => sinef <= 8099;
 when 1123 => sinef <= 8097;
 when 1124 => sinef <= 8095;
 when 1125 => sinef <= 8093;
 when 1126 => sinef <= 8091;
 when 1127 => sinef <= 8089;
 when 1128 => sinef <= 8087;
 when 1129 => sinef <= 8085;
 when 1130 => sinef <= 8083;
 when 1131 => sinef <= 8081;
 when 1132 => sinef <= 8079;
 when 1133 => sinef <= 8077;
 when 1134 => sinef <= 8075;
 when 1135 => sinef <= 8073;
 when 1136 => sinef <= 8070;
 when 1137 => sinef <= 8068;
 when 1138 => sinef <= 8066;
 when 1139 => sinef <= 8064;
 when 1140 => sinef <= 8062;
 when 1141 => sinef <= 8059;
 when 1142 => sinef <= 8057;
 when 1143 => sinef <= 8055;
 when 1144 => sinef <= 8053;
 when 1145 => sinef <= 8050;
 when 1146 => sinef <= 8048;
 when 1147 => sinef <= 8046;
 when 1148 => sinef <= 8043;
 when 1149 => sinef <= 8041;
 when 1150 => sinef <= 8038;
 when 1151 => sinef <= 8036;
 when 1152 => sinef <= 8034;
 when 1153 => sinef <= 8031;
 when 1154 => sinef <= 8029;
 when 1155 => sinef <= 8026;
 when 1156 => sinef <= 8024;
 when 1157 => sinef <= 8021;
 when 1158 => sinef <= 8019;
 when 1159 => sinef <= 8016;
 when 1160 => sinef <= 8013;
 when 1161 => sinef <= 8011;
 when 1162 => sinef <= 8008;
 when 1163 => sinef <= 8006;
 when 1164 => sinef <= 8003;
 when 1165 => sinef <= 8000;
 when 1166 => sinef <= 7997;
 when 1167 => sinef <= 7995;
 when 1168 => sinef <= 7992;
 when 1169 => sinef <= 7989;
 when 1170 => sinef <= 7986;
 when 1171 => sinef <= 7984;
 when 1172 => sinef <= 7981;
 when 1173 => sinef <= 7978;
 when 1174 => sinef <= 7975;
 when 1175 => sinef <= 7972;
 when 1176 => sinef <= 7969;
 when 1177 => sinef <= 7966;
 when 1178 => sinef <= 7964;
 when 1179 => sinef <= 7961;
 when 1180 => sinef <= 7958;
 when 1181 => sinef <= 7955;
 when 1182 => sinef <= 7952;
 when 1183 => sinef <= 7949;
 when 1184 => sinef <= 7946;
 when 1185 => sinef <= 7942;
 when 1186 => sinef <= 7939;
 when 1187 => sinef <= 7936;
 when 1188 => sinef <= 7933;
 when 1189 => sinef <= 7930;
 when 1190 => sinef <= 7927;
 when 1191 => sinef <= 7924;
 when 1192 => sinef <= 7921;
 when 1193 => sinef <= 7917;
 when 1194 => sinef <= 7914;
 when 1195 => sinef <= 7911;
 when 1196 => sinef <= 7908;
 when 1197 => sinef <= 7904;
 when 1198 => sinef <= 7901;
 when 1199 => sinef <= 7898;
 when 1200 => sinef <= 7894;
 when 1201 => sinef <= 7891;
 when 1202 => sinef <= 7888;
 when 1203 => sinef <= 7884;
 when 1204 => sinef <= 7881;
 when 1205 => sinef <= 7877;
 when 1206 => sinef <= 7874;
 when 1207 => sinef <= 7870;
 when 1208 => sinef <= 7867;
 when 1209 => sinef <= 7863;
 when 1210 => sinef <= 7860;
 when 1211 => sinef <= 7856;
 when 1212 => sinef <= 7853;
 when 1213 => sinef <= 7849;
 when 1214 => sinef <= 7846;
 when 1215 => sinef <= 7842;
 when 1216 => sinef <= 7838;
 when 1217 => sinef <= 7835;
 when 1218 => sinef <= 7831;
 when 1219 => sinef <= 7827;
 when 1220 => sinef <= 7824;
 when 1221 => sinef <= 7820;
 when 1222 => sinef <= 7816;
 when 1223 => sinef <= 7812;
 when 1224 => sinef <= 7809;
 when 1225 => sinef <= 7805;
 when 1226 => sinef <= 7801;
 when 1227 => sinef <= 7797;
 when 1228 => sinef <= 7793;
 when 1229 => sinef <= 7789;
 when 1230 => sinef <= 7785;
 when 1231 => sinef <= 7782;
 when 1232 => sinef <= 7778;
 when 1233 => sinef <= 7774;
 when 1234 => sinef <= 7770;
 when 1235 => sinef <= 7766;
 when 1236 => sinef <= 7762;
 when 1237 => sinef <= 7758;
 when 1238 => sinef <= 7754;
 when 1239 => sinef <= 7750;
 when 1240 => sinef <= 7745;
 when 1241 => sinef <= 7741;
 when 1242 => sinef <= 7737;
 when 1243 => sinef <= 7733;
 when 1244 => sinef <= 7729;
 when 1245 => sinef <= 7725;
 when 1246 => sinef <= 7721;
 when 1247 => sinef <= 7716;
 when 1248 => sinef <= 7712;
 when 1249 => sinef <= 7708;
 when 1250 => sinef <= 7704;
 when 1251 => sinef <= 7699;
 when 1252 => sinef <= 7695;
 when 1253 => sinef <= 7691;
 when 1254 => sinef <= 7686;
 when 1255 => sinef <= 7682;
 when 1256 => sinef <= 7678;
 when 1257 => sinef <= 7673;
 when 1258 => sinef <= 7669;
 when 1259 => sinef <= 7665;
 when 1260 => sinef <= 7660;
 when 1261 => sinef <= 7656;
 when 1262 => sinef <= 7651;
 when 1263 => sinef <= 7647;
 when 1264 => sinef <= 7642;
 when 1265 => sinef <= 7638;
 when 1266 => sinef <= 7633;
 when 1267 => sinef <= 7628;
 when 1268 => sinef <= 7624;
 when 1269 => sinef <= 7619;
 when 1270 => sinef <= 7615;
 when 1271 => sinef <= 7610;
 when 1272 => sinef <= 7605;
 when 1273 => sinef <= 7601;
 when 1274 => sinef <= 7596;
 when 1275 => sinef <= 7591;
 when 1276 => sinef <= 7587;
 when 1277 => sinef <= 7582;
 when 1278 => sinef <= 7577;
 when 1279 => sinef <= 7572;
 when 1280 => sinef <= 7567;
 when 1281 => sinef <= 7563;
 when 1282 => sinef <= 7558;
 when 1283 => sinef <= 7553;
 when 1284 => sinef <= 7548;
 when 1285 => sinef <= 7543;
 when 1286 => sinef <= 7538;
 when 1287 => sinef <= 7533;
 when 1288 => sinef <= 7528;
 when 1289 => sinef <= 7524;
 when 1290 => sinef <= 7519;
 when 1291 => sinef <= 7514;
 when 1292 => sinef <= 7509;
 when 1293 => sinef <= 7503;
 when 1294 => sinef <= 7498;
 when 1295 => sinef <= 7493;
 when 1296 => sinef <= 7488;
 when 1297 => sinef <= 7483;
 when 1298 => sinef <= 7478;
 when 1299 => sinef <= 7473;
 when 1300 => sinef <= 7468;
 when 1301 => sinef <= 7463;
 when 1302 => sinef <= 7457;
 when 1303 => sinef <= 7452;
 when 1304 => sinef <= 7447;
 when 1305 => sinef <= 7442;
 when 1306 => sinef <= 7436;
 when 1307 => sinef <= 7431;
 when 1308 => sinef <= 7426;
 when 1309 => sinef <= 7421;
 when 1310 => sinef <= 7415;
 when 1311 => sinef <= 7410;
 when 1312 => sinef <= 7405;
 when 1313 => sinef <= 7399;
 when 1314 => sinef <= 7394;
 when 1315 => sinef <= 7388;
 when 1316 => sinef <= 7383;
 when 1317 => sinef <= 7377;
 when 1318 => sinef <= 7372;
 when 1319 => sinef <= 7367;
 when 1320 => sinef <= 7361;
 when 1321 => sinef <= 7356;
 when 1322 => sinef <= 7350;
 when 1323 => sinef <= 7344;
 when 1324 => sinef <= 7339;
 when 1325 => sinef <= 7333;
 when 1326 => sinef <= 7328;
 when 1327 => sinef <= 7322;
 when 1328 => sinef <= 7316;
 when 1329 => sinef <= 7311;
 when 1330 => sinef <= 7305;
 when 1331 => sinef <= 7299;
 when 1332 => sinef <= 7294;
 when 1333 => sinef <= 7288;
 when 1334 => sinef <= 7282;
 when 1335 => sinef <= 7276;
 when 1336 => sinef <= 7271;
 when 1337 => sinef <= 7265;
 when 1338 => sinef <= 7259;
 when 1339 => sinef <= 7253;
 when 1340 => sinef <= 7247;
 when 1341 => sinef <= 7242;
 when 1342 => sinef <= 7236;
 when 1343 => sinef <= 7230;
 when 1344 => sinef <= 7224;
 when 1345 => sinef <= 7218;
 when 1346 => sinef <= 7212;
 when 1347 => sinef <= 7206;
 when 1348 => sinef <= 7200;
 when 1349 => sinef <= 7194;
 when 1350 => sinef <= 7188;
 when 1351 => sinef <= 7182;
 when 1352 => sinef <= 7176;
 when 1353 => sinef <= 7170;
 when 1354 => sinef <= 7164;
 when 1355 => sinef <= 7158;
 when 1356 => sinef <= 7152;
 when 1357 => sinef <= 7145;
 when 1358 => sinef <= 7139;
 when 1359 => sinef <= 7133;
 when 1360 => sinef <= 7127;
 when 1361 => sinef <= 7121;
 when 1362 => sinef <= 7114;
 when 1363 => sinef <= 7108;
 when 1364 => sinef <= 7102;
 when 1365 => sinef <= 7096;
 when 1366 => sinef <= 7089;
 when 1367 => sinef <= 7083;
 when 1368 => sinef <= 7077;
 when 1369 => sinef <= 7070;
 when 1370 => sinef <= 7064;
 when 1371 => sinef <= 7058;
 when 1372 => sinef <= 7051;
 when 1373 => sinef <= 7045;
 when 1374 => sinef <= 7039;
 when 1375 => sinef <= 7032;
 when 1376 => sinef <= 7026;
 when 1377 => sinef <= 7019;
 when 1378 => sinef <= 7013;
 when 1379 => sinef <= 7006;
 when 1380 => sinef <= 7000;
 when 1381 => sinef <= 6993;
 when 1382 => sinef <= 6987;
 when 1383 => sinef <= 6980;
 when 1384 => sinef <= 6973;
 when 1385 => sinef <= 6967;
 when 1386 => sinef <= 6960;
 when 1387 => sinef <= 6954;
 when 1388 => sinef <= 6947;
 when 1389 => sinef <= 6940;
 when 1390 => sinef <= 6934;
 when 1391 => sinef <= 6927;
 when 1392 => sinef <= 6920;
 when 1393 => sinef <= 6913;
 when 1394 => sinef <= 6907;
 when 1395 => sinef <= 6900;
 when 1396 => sinef <= 6893;
 when 1397 => sinef <= 6886;
 when 1398 => sinef <= 6880;
 when 1399 => sinef <= 6873;
 when 1400 => sinef <= 6866;
 when 1401 => sinef <= 6859;
 when 1402 => sinef <= 6852;
 when 1403 => sinef <= 6845;
 when 1404 => sinef <= 6838;
 when 1405 => sinef <= 6831;
 when 1406 => sinef <= 6824;
 when 1407 => sinef <= 6818;
 when 1408 => sinef <= 6811;
 when 1409 => sinef <= 6804;
 when 1410 => sinef <= 6797;
 when 1411 => sinef <= 6790;
 when 1412 => sinef <= 6783;
 when 1413 => sinef <= 6775;
 when 1414 => sinef <= 6768;
 when 1415 => sinef <= 6761;
 when 1416 => sinef <= 6754;
 when 1417 => sinef <= 6747;
 when 1418 => sinef <= 6740;
 when 1419 => sinef <= 6733;
 when 1420 => sinef <= 6726;
 when 1421 => sinef <= 6718;
 when 1422 => sinef <= 6711;
 when 1423 => sinef <= 6704;
 when 1424 => sinef <= 6697;
 when 1425 => sinef <= 6690;
 when 1426 => sinef <= 6682;
 when 1427 => sinef <= 6675;
 when 1428 => sinef <= 6668;
 when 1429 => sinef <= 6660;
 when 1430 => sinef <= 6653;
 when 1431 => sinef <= 6646;
 when 1432 => sinef <= 6638;
 when 1433 => sinef <= 6631;
 when 1434 => sinef <= 6624;
 when 1435 => sinef <= 6616;
 when 1436 => sinef <= 6609;
 when 1437 => sinef <= 6601;
 when 1438 => sinef <= 6594;
 when 1439 => sinef <= 6587;
 when 1440 => sinef <= 6579;
 when 1441 => sinef <= 6572;
 when 1442 => sinef <= 6564;
 when 1443 => sinef <= 6557;
 when 1444 => sinef <= 6549;
 when 1445 => sinef <= 6541;
 when 1446 => sinef <= 6534;
 when 1447 => sinef <= 6526;
 when 1448 => sinef <= 6519;
 when 1449 => sinef <= 6511;
 when 1450 => sinef <= 6503;
 when 1451 => sinef <= 6496;
 when 1452 => sinef <= 6488;
 when 1453 => sinef <= 6480;
 when 1454 => sinef <= 6473;
 when 1455 => sinef <= 6465;
 when 1456 => sinef <= 6457;
 when 1457 => sinef <= 6450;
 when 1458 => sinef <= 6442;
 when 1459 => sinef <= 6434;
 when 1460 => sinef <= 6426;
 when 1461 => sinef <= 6419;
 when 1462 => sinef <= 6411;
 when 1463 => sinef <= 6403;
 when 1464 => sinef <= 6395;
 when 1465 => sinef <= 6387;
 when 1466 => sinef <= 6379;
 when 1467 => sinef <= 6371;
 when 1468 => sinef <= 6363;
 when 1469 => sinef <= 6356;
 when 1470 => sinef <= 6348;
 when 1471 => sinef <= 6340;
 when 1472 => sinef <= 6332;
 when 1473 => sinef <= 6324;
 when 1474 => sinef <= 6316;
 when 1475 => sinef <= 6308;
 when 1476 => sinef <= 6300;
 when 1477 => sinef <= 6292;
 when 1478 => sinef <= 6284;
 when 1479 => sinef <= 6276;
 when 1480 => sinef <= 6267;
 when 1481 => sinef <= 6259;
 when 1482 => sinef <= 6251;
 when 1483 => sinef <= 6243;
 when 1484 => sinef <= 6235;
 when 1485 => sinef <= 6227;
 when 1486 => sinef <= 6219;
 when 1487 => sinef <= 6210;
 when 1488 => sinef <= 6202;
 when 1489 => sinef <= 6194;
 when 1490 => sinef <= 6186;
 when 1491 => sinef <= 6178;
 when 1492 => sinef <= 6169;
 when 1493 => sinef <= 6161;
 when 1494 => sinef <= 6153;
 when 1495 => sinef <= 6144;
 when 1496 => sinef <= 6136;
 when 1497 => sinef <= 6128;
 when 1498 => sinef <= 6120;
 when 1499 => sinef <= 6111;
 when 1500 => sinef <= 6103;
 when 1501 => sinef <= 6094;
 when 1502 => sinef <= 6086;
 when 1503 => sinef <= 6078;
 when 1504 => sinef <= 6069;
 when 1505 => sinef <= 6061;
 when 1506 => sinef <= 6052;
 when 1507 => sinef <= 6044;
 when 1508 => sinef <= 6035;
 when 1509 => sinef <= 6027;
 when 1510 => sinef <= 6018;
 when 1511 => sinef <= 6010;
 when 1512 => sinef <= 6001;
 when 1513 => sinef <= 5993;
 when 1514 => sinef <= 5984;
 when 1515 => sinef <= 5975;
 when 1516 => sinef <= 5967;
 when 1517 => sinef <= 5958;
 when 1518 => sinef <= 5950;
 when 1519 => sinef <= 5941;
 when 1520 => sinef <= 5932;
 when 1521 => sinef <= 5924;
 when 1522 => sinef <= 5915;
 when 1523 => sinef <= 5906;
 when 1524 => sinef <= 5898;
 when 1525 => sinef <= 5889;
 when 1526 => sinef <= 5880;
 when 1527 => sinef <= 5871;
 when 1528 => sinef <= 5863;
 when 1529 => sinef <= 5854;
 when 1530 => sinef <= 5845;
 when 1531 => sinef <= 5836;
 when 1532 => sinef <= 5827;
 when 1533 => sinef <= 5819;
 when 1534 => sinef <= 5810;
 when 1535 => sinef <= 5801;
 when 1536 => sinef <= 5792;
 when 1537 => sinef <= 5783;
 when 1538 => sinef <= 5774;
 when 1539 => sinef <= 5765;
 when 1540 => sinef <= 5756;
 when 1541 => sinef <= 5747;
 when 1542 => sinef <= 5738;
 when 1543 => sinef <= 5729;
 when 1544 => sinef <= 5720;
 when 1545 => sinef <= 5711;
 when 1546 => sinef <= 5702;
 when 1547 => sinef <= 5693;
 when 1548 => sinef <= 5684;
 when 1549 => sinef <= 5675;
 when 1550 => sinef <= 5666;
 when 1551 => sinef <= 5657;
 when 1552 => sinef <= 5648;
 when 1553 => sinef <= 5639;
 when 1554 => sinef <= 5630;
 when 1555 => sinef <= 5621;
 when 1556 => sinef <= 5612;
 when 1557 => sinef <= 5602;
 when 1558 => sinef <= 5593;
 when 1559 => sinef <= 5584;
 when 1560 => sinef <= 5575;
 when 1561 => sinef <= 5566;
 when 1562 => sinef <= 5556;
 when 1563 => sinef <= 5547;
 when 1564 => sinef <= 5538;
 when 1565 => sinef <= 5529;
 when 1566 => sinef <= 5519;
 when 1567 => sinef <= 5510;
 when 1568 => sinef <= 5501;
 when 1569 => sinef <= 5491;
 when 1570 => sinef <= 5482;
 when 1571 => sinef <= 5473;
 when 1572 => sinef <= 5463;
 when 1573 => sinef <= 5454;
 when 1574 => sinef <= 5445;
 when 1575 => sinef <= 5435;
 when 1576 => sinef <= 5426;
 when 1577 => sinef <= 5416;
 when 1578 => sinef <= 5407;
 when 1579 => sinef <= 5398;
 when 1580 => sinef <= 5388;
 when 1581 => sinef <= 5379;
 when 1582 => sinef <= 5369;
 when 1583 => sinef <= 5360;
 when 1584 => sinef <= 5350;
 when 1585 => sinef <= 5341;
 when 1586 => sinef <= 5331;
 when 1587 => sinef <= 5322;
 when 1588 => sinef <= 5312;
 when 1589 => sinef <= 5302;
 when 1590 => sinef <= 5293;
 when 1591 => sinef <= 5283;
 when 1592 => sinef <= 5274;
 when 1593 => sinef <= 5264;
 when 1594 => sinef <= 5254;
 when 1595 => sinef <= 5245;
 when 1596 => sinef <= 5235;
 when 1597 => sinef <= 5225;
 when 1598 => sinef <= 5216;
 when 1599 => sinef <= 5206;
 when 1600 => sinef <= 5196;
 when 1601 => sinef <= 5187;
 when 1602 => sinef <= 5177;
 when 1603 => sinef <= 5167;
 when 1604 => sinef <= 5157;
 when 1605 => sinef <= 5148;
 when 1606 => sinef <= 5138;
 when 1607 => sinef <= 5128;
 when 1608 => sinef <= 5118;
 when 1609 => sinef <= 5108;
 when 1610 => sinef <= 5099;
 when 1611 => sinef <= 5089;
 when 1612 => sinef <= 5079;
 when 1613 => sinef <= 5069;
 when 1614 => sinef <= 5059;
 when 1615 => sinef <= 5049;
 when 1616 => sinef <= 5039;
 when 1617 => sinef <= 5029;
 when 1618 => sinef <= 5020;
 when 1619 => sinef <= 5010;
 when 1620 => sinef <= 5000;
 when 1621 => sinef <= 4990;
 when 1622 => sinef <= 4980;
 when 1623 => sinef <= 4970;
 when 1624 => sinef <= 4960;
 when 1625 => sinef <= 4950;
 when 1626 => sinef <= 4940;
 when 1627 => sinef <= 4930;
 when 1628 => sinef <= 4920;
 when 1629 => sinef <= 4910;
 when 1630 => sinef <= 4900;
 when 1631 => sinef <= 4889;
 when 1632 => sinef <= 4879;
 when 1633 => sinef <= 4869;
 when 1634 => sinef <= 4859;
 when 1635 => sinef <= 4849;
 when 1636 => sinef <= 4839;
 when 1637 => sinef <= 4829;
 when 1638 => sinef <= 4819;
 when 1639 => sinef <= 4808;
 when 1640 => sinef <= 4798;
 when 1641 => sinef <= 4788;
 when 1642 => sinef <= 4778;
 when 1643 => sinef <= 4768;
 when 1644 => sinef <= 4757;
 when 1645 => sinef <= 4747;
 when 1646 => sinef <= 4737;
 when 1647 => sinef <= 4727;
 when 1648 => sinef <= 4716;
 when 1649 => sinef <= 4706;
 when 1650 => sinef <= 4696;
 when 1651 => sinef <= 4686;
 when 1652 => sinef <= 4675;
 when 1653 => sinef <= 4665;
 when 1654 => sinef <= 4655;
 when 1655 => sinef <= 4644;
 when 1656 => sinef <= 4634;
 when 1657 => sinef <= 4624;
 when 1658 => sinef <= 4613;
 when 1659 => sinef <= 4603;
 when 1660 => sinef <= 4592;
 when 1661 => sinef <= 4582;
 when 1662 => sinef <= 4572;
 when 1663 => sinef <= 4561;
 when 1664 => sinef <= 4551;
 when 1665 => sinef <= 4540;
 when 1666 => sinef <= 4530;
 when 1667 => sinef <= 4519;
 when 1668 => sinef <= 4509;
 when 1669 => sinef <= 4498;
 when 1670 => sinef <= 4488;
 when 1671 => sinef <= 4477;
 when 1672 => sinef <= 4467;
 when 1673 => sinef <= 4456;
 when 1674 => sinef <= 4446;
 when 1675 => sinef <= 4435;
 when 1676 => sinef <= 4425;
 when 1677 => sinef <= 4414;
 when 1678 => sinef <= 4403;
 when 1679 => sinef <= 4393;
 when 1680 => sinef <= 4382;
 when 1681 => sinef <= 4372;
 when 1682 => sinef <= 4361;
 when 1683 => sinef <= 4350;
 when 1684 => sinef <= 4340;
 when 1685 => sinef <= 4329;
 when 1686 => sinef <= 4318;
 when 1687 => sinef <= 4308;
 when 1688 => sinef <= 4297;
 when 1689 => sinef <= 4286;
 when 1690 => sinef <= 4275;
 when 1691 => sinef <= 4265;
 when 1692 => sinef <= 4254;
 when 1693 => sinef <= 4243;
 when 1694 => sinef <= 4233;
 when 1695 => sinef <= 4222;
 when 1696 => sinef <= 4211;
 when 1697 => sinef <= 4200;
 when 1698 => sinef <= 4189;
 when 1699 => sinef <= 4179;
 when 1700 => sinef <= 4168;
 when 1701 => sinef <= 4157;
 when 1702 => sinef <= 4146;
 when 1703 => sinef <= 4135;
 when 1704 => sinef <= 4124;
 when 1705 => sinef <= 4114;
 when 1706 => sinef <= 4103;
 when 1707 => sinef <= 4092;
 when 1708 => sinef <= 4081;
 when 1709 => sinef <= 4070;
 when 1710 => sinef <= 4059;
 when 1711 => sinef <= 4048;
 when 1712 => sinef <= 4037;
 when 1713 => sinef <= 4026;
 when 1714 => sinef <= 4015;
 when 1715 => sinef <= 4004;
 when 1716 => sinef <= 3994;
 when 1717 => sinef <= 3983;
 when 1718 => sinef <= 3972;
 when 1719 => sinef <= 3961;
 when 1720 => sinef <= 3950;
 when 1721 => sinef <= 3939;
 when 1722 => sinef <= 3928;
 when 1723 => sinef <= 3917;
 when 1724 => sinef <= 3905;
 when 1725 => sinef <= 3894;
 when 1726 => sinef <= 3883;
 when 1727 => sinef <= 3872;
 when 1728 => sinef <= 3861;
 when 1729 => sinef <= 3850;
 when 1730 => sinef <= 3839;
 when 1731 => sinef <= 3828;
 when 1732 => sinef <= 3817;
 when 1733 => sinef <= 3806;
 when 1734 => sinef <= 3795;
 when 1735 => sinef <= 3783;
 when 1736 => sinef <= 3772;
 when 1737 => sinef <= 3761;
 when 1738 => sinef <= 3750;
 when 1739 => sinef <= 3739;
 when 1740 => sinef <= 3728;
 when 1741 => sinef <= 3716;
 when 1742 => sinef <= 3705;
 when 1743 => sinef <= 3694;
 when 1744 => sinef <= 3683;
 when 1745 => sinef <= 3672;
 when 1746 => sinef <= 3660;
 when 1747 => sinef <= 3649;
 when 1748 => sinef <= 3638;
 when 1749 => sinef <= 3627;
 when 1750 => sinef <= 3615;
 when 1751 => sinef <= 3604;
 when 1752 => sinef <= 3593;
 when 1753 => sinef <= 3581;
 when 1754 => sinef <= 3570;
 when 1755 => sinef <= 3559;
 when 1756 => sinef <= 3547;
 when 1757 => sinef <= 3536;
 when 1758 => sinef <= 3525;
 when 1759 => sinef <= 3513;
 when 1760 => sinef <= 3502;
 when 1761 => sinef <= 3491;
 when 1762 => sinef <= 3479;
 when 1763 => sinef <= 3468;
 when 1764 => sinef <= 3457;
 when 1765 => sinef <= 3445;
 when 1766 => sinef <= 3434;
 when 1767 => sinef <= 3422;
 when 1768 => sinef <= 3411;
 when 1769 => sinef <= 3400;
 when 1770 => sinef <= 3388;
 when 1771 => sinef <= 3377;
 when 1772 => sinef <= 3365;
 when 1773 => sinef <= 3354;
 when 1774 => sinef <= 3342;
 when 1775 => sinef <= 3331;
 when 1776 => sinef <= 3319;
 when 1777 => sinef <= 3308;
 when 1778 => sinef <= 3296;
 when 1779 => sinef <= 3285;
 when 1780 => sinef <= 3273;
 when 1781 => sinef <= 3262;
 when 1782 => sinef <= 3250;
 when 1783 => sinef <= 3239;
 when 1784 => sinef <= 3227;
 when 1785 => sinef <= 3216;
 when 1786 => sinef <= 3204;
 when 1787 => sinef <= 3193;
 when 1788 => sinef <= 3181;
 when 1789 => sinef <= 3169;
 when 1790 => sinef <= 3158;
 when 1791 => sinef <= 3146;
 when 1792 => sinef <= 3135;
 when 1793 => sinef <= 3123;
 when 1794 => sinef <= 3111;
 when 1795 => sinef <= 3100;
 when 1796 => sinef <= 3088;
 when 1797 => sinef <= 3076;
 when 1798 => sinef <= 3065;
 when 1799 => sinef <= 3053;
 when 1800 => sinef <= 3041;
 when 1801 => sinef <= 3030;
 when 1802 => sinef <= 3018;
 when 1803 => sinef <= 3006;
 when 1804 => sinef <= 2995;
 when 1805 => sinef <= 2983;
 when 1806 => sinef <= 2971;
 when 1807 => sinef <= 2960;
 when 1808 => sinef <= 2948;
 when 1809 => sinef <= 2936;
 when 1810 => sinef <= 2924;
 when 1811 => sinef <= 2913;
 when 1812 => sinef <= 2901;
 when 1813 => sinef <= 2889;
 when 1814 => sinef <= 2877;
 when 1815 => sinef <= 2866;
 when 1816 => sinef <= 2854;
 when 1817 => sinef <= 2842;
 when 1818 => sinef <= 2830;
 when 1819 => sinef <= 2819;
 when 1820 => sinef <= 2807;
 when 1821 => sinef <= 2795;
 when 1822 => sinef <= 2783;
 when 1823 => sinef <= 2771;
 when 1824 => sinef <= 2759;
 when 1825 => sinef <= 2748;
 when 1826 => sinef <= 2736;
 when 1827 => sinef <= 2724;
 when 1828 => sinef <= 2712;
 when 1829 => sinef <= 2700;
 when 1830 => sinef <= 2688;
 when 1831 => sinef <= 2676;
 when 1832 => sinef <= 2665;
 when 1833 => sinef <= 2653;
 when 1834 => sinef <= 2641;
 when 1835 => sinef <= 2629;
 when 1836 => sinef <= 2617;
 when 1837 => sinef <= 2605;
 when 1838 => sinef <= 2593;
 when 1839 => sinef <= 2581;
 when 1840 => sinef <= 2569;
 when 1841 => sinef <= 2557;
 when 1842 => sinef <= 2545;
 when 1843 => sinef <= 2534;
 when 1844 => sinef <= 2522;
 when 1845 => sinef <= 2510;
 when 1846 => sinef <= 2498;
 when 1847 => sinef <= 2486;
 when 1848 => sinef <= 2474;
 when 1849 => sinef <= 2462;
 when 1850 => sinef <= 2450;
 when 1851 => sinef <= 2438;
 when 1852 => sinef <= 2426;
 when 1853 => sinef <= 2414;
 when 1854 => sinef <= 2402;
 when 1855 => sinef <= 2390;
 when 1856 => sinef <= 2378;
 when 1857 => sinef <= 2366;
 when 1858 => sinef <= 2354;
 when 1859 => sinef <= 2342;
 when 1860 => sinef <= 2330;
 when 1861 => sinef <= 2318;
 when 1862 => sinef <= 2305;
 when 1863 => sinef <= 2293;
 when 1864 => sinef <= 2281;
 when 1865 => sinef <= 2269;
 when 1866 => sinef <= 2257;
 when 1867 => sinef <= 2245;
 when 1868 => sinef <= 2233;
 when 1869 => sinef <= 2221;
 when 1870 => sinef <= 2209;
 when 1871 => sinef <= 2197;
 when 1872 => sinef <= 2185;
 when 1873 => sinef <= 2173;
 when 1874 => sinef <= 2160;
 when 1875 => sinef <= 2148;
 when 1876 => sinef <= 2136;
 when 1877 => sinef <= 2124;
 when 1878 => sinef <= 2112;
 when 1879 => sinef <= 2100;
 when 1880 => sinef <= 2088;
 when 1881 => sinef <= 2075;
 when 1882 => sinef <= 2063;
 when 1883 => sinef <= 2051;
 when 1884 => sinef <= 2039;
 when 1885 => sinef <= 2027;
 when 1886 => sinef <= 2015;
 when 1887 => sinef <= 2002;
 when 1888 => sinef <= 1990;
 when 1889 => sinef <= 1978;
 when 1890 => sinef <= 1966;
 when 1891 => sinef <= 1954;
 when 1892 => sinef <= 1941;
 when 1893 => sinef <= 1929;
 when 1894 => sinef <= 1917;
 when 1895 => sinef <= 1905;
 when 1896 => sinef <= 1893;
 when 1897 => sinef <= 1880;
 when 1898 => sinef <= 1868;
 when 1899 => sinef <= 1856;
 when 1900 => sinef <= 1844;
 when 1901 => sinef <= 1831;
 when 1902 => sinef <= 1819;
 when 1903 => sinef <= 1807;
 when 1904 => sinef <= 1795;
 when 1905 => sinef <= 1782;
 when 1906 => sinef <= 1770;
 when 1907 => sinef <= 1758;
 when 1908 => sinef <= 1746;
 when 1909 => sinef <= 1733;
 when 1910 => sinef <= 1721;
 when 1911 => sinef <= 1709;
 when 1912 => sinef <= 1696;
 when 1913 => sinef <= 1684;
 when 1914 => sinef <= 1672;
 when 1915 => sinef <= 1660;
 when 1916 => sinef <= 1647;
 when 1917 => sinef <= 1635;
 when 1918 => sinef <= 1623;
 when 1919 => sinef <= 1610;
 when 1920 => sinef <= 1598;
 when 1921 => sinef <= 1586;
 when 1922 => sinef <= 1573;
 when 1923 => sinef <= 1561;
 when 1924 => sinef <= 1549;
 when 1925 => sinef <= 1536;
 when 1926 => sinef <= 1524;
 when 1927 => sinef <= 1512;
 when 1928 => sinef <= 1499;
 when 1929 => sinef <= 1487;
 when 1930 => sinef <= 1475;
 when 1931 => sinef <= 1462;
 when 1932 => sinef <= 1450;
 when 1933 => sinef <= 1437;
 when 1934 => sinef <= 1425;
 when 1935 => sinef <= 1413;
 when 1936 => sinef <= 1400;
 when 1937 => sinef <= 1388;
 when 1938 => sinef <= 1376;
 when 1939 => sinef <= 1363;
 when 1940 => sinef <= 1351;
 when 1941 => sinef <= 1338;
 when 1942 => sinef <= 1326;
 when 1943 => sinef <= 1314;
 when 1944 => sinef <= 1301;
 when 1945 => sinef <= 1289;
 when 1946 => sinef <= 1276;
 when 1947 => sinef <= 1264;
 when 1948 => sinef <= 1252;
 when 1949 => sinef <= 1239;
 when 1950 => sinef <= 1227;
 when 1951 => sinef <= 1214;
 when 1952 => sinef <= 1202;
 when 1953 => sinef <= 1189;
 when 1954 => sinef <= 1177;
 when 1955 => sinef <= 1165;
 when 1956 => sinef <= 1152;
 when 1957 => sinef <= 1140;
 when 1958 => sinef <= 1127;
 when 1959 => sinef <= 1115;
 when 1960 => sinef <= 1102;
 when 1961 => sinef <= 1090;
 when 1962 => sinef <= 1077;
 when 1963 => sinef <= 1065;
 when 1964 => sinef <= 1053;
 when 1965 => sinef <= 1040;
 when 1966 => sinef <= 1028;
 when 1967 => sinef <= 1015;
 when 1968 => sinef <= 1003;
 when 1969 => sinef <= 990;
 when 1970 => sinef <= 978;
 when 1971 => sinef <= 965;
 when 1972 => sinef <= 953;
 when 1973 => sinef <= 940;
 when 1974 => sinef <= 928;
 when 1975 => sinef <= 915;
 when 1976 => sinef <= 903;
 when 1977 => sinef <= 890;
 when 1978 => sinef <= 878;
 when 1979 => sinef <= 865;
 when 1980 => sinef <= 853;
 when 1981 => sinef <= 840;
 when 1982 => sinef <= 828;
 when 1983 => sinef <= 815;
 when 1984 => sinef <= 803;
 when 1985 => sinef <= 790;
 when 1986 => sinef <= 778;
 when 1987 => sinef <= 765;
 when 1988 => sinef <= 753;
 when 1989 => sinef <= 740;
 when 1990 => sinef <= 728;
 when 1991 => sinef <= 715;
 when 1992 => sinef <= 703;
 when 1993 => sinef <= 690;
 when 1994 => sinef <= 678;
 when 1995 => sinef <= 665;
 when 1996 => sinef <= 653;
 when 1997 => sinef <= 640;
 when 1998 => sinef <= 628;
 when 1999 => sinef <= 615;
 when 2000 => sinef <= 603;
 when 2001 => sinef <= 590;
 when 2002 => sinef <= 578;
 when 2003 => sinef <= 565;
 when 2004 => sinef <= 552;
 when 2005 => sinef <= 540;
 when 2006 => sinef <= 527;
 when 2007 => sinef <= 515;
 when 2008 => sinef <= 502;
 when 2009 => sinef <= 490;
 when 2010 => sinef <= 477;
 when 2011 => sinef <= 465;
 when 2012 => sinef <= 452;
 when 2013 => sinef <= 440;
 when 2014 => sinef <= 427;
 when 2015 => sinef <= 414;
 when 2016 => sinef <= 402;
 when 2017 => sinef <= 389;
 when 2018 => sinef <= 377;
 when 2019 => sinef <= 364;
 when 2020 => sinef <= 352;
 when 2021 => sinef <= 339;
 when 2022 => sinef <= 327;
 when 2023 => sinef <= 314;
 when 2024 => sinef <= 301;
 when 2025 => sinef <= 289;
 when 2026 => sinef <= 276;
 when 2027 => sinef <= 264;
 when 2028 => sinef <= 251;
 when 2029 => sinef <= 239;
 when 2030 => sinef <= 226;
 when 2031 => sinef <= 214;
 when 2032 => sinef <= 201;
 when 2033 => sinef <= 188;
 when 2034 => sinef <= 176;
 when 2035 => sinef <= 163;
 when 2036 => sinef <= 151;
 when 2037 => sinef <= 138;
 when 2038 => sinef <= 126;
 when 2039 => sinef <= 113;
 when 2040 => sinef <= 101;
 when 2041 => sinef <= 88;
 when 2042 => sinef <= 75;
 when 2043 => sinef <= 63;
 when 2044 => sinef <= 50;
 when 2045 => sinef <= 38;
 when 2046 => sinef <= 25;
 when 2047 => sinef <= 13;
 when 2048 => sinef <= 0;
 when 2049 => sinef <= -13;
 when 2050 => sinef <= -25;
 when 2051 => sinef <= -38;
 when 2052 => sinef <= -50;
 when 2053 => sinef <= -63;
 when 2054 => sinef <= -75;
 when 2055 => sinef <= -88;
 when 2056 => sinef <= -101;
 when 2057 => sinef <= -113;
 when 2058 => sinef <= -126;
 when 2059 => sinef <= -138;
 when 2060 => sinef <= -151;
 when 2061 => sinef <= -163;
 when 2062 => sinef <= -176;
 when 2063 => sinef <= -188;
 when 2064 => sinef <= -201;
 when 2065 => sinef <= -214;
 when 2066 => sinef <= -226;
 when 2067 => sinef <= -239;
 when 2068 => sinef <= -251;
 when 2069 => sinef <= -264;
 when 2070 => sinef <= -276;
 when 2071 => sinef <= -289;
 when 2072 => sinef <= -301;
 when 2073 => sinef <= -314;
 when 2074 => sinef <= -327;
 when 2075 => sinef <= -339;
 when 2076 => sinef <= -352;
 when 2077 => sinef <= -364;
 when 2078 => sinef <= -377;
 when 2079 => sinef <= -389;
 when 2080 => sinef <= -402;
 when 2081 => sinef <= -414;
 when 2082 => sinef <= -427;
 when 2083 => sinef <= -440;
 when 2084 => sinef <= -452;
 when 2085 => sinef <= -465;
 when 2086 => sinef <= -477;
 when 2087 => sinef <= -490;
 when 2088 => sinef <= -502;
 when 2089 => sinef <= -515;
 when 2090 => sinef <= -527;
 when 2091 => sinef <= -540;
 when 2092 => sinef <= -552;
 when 2093 => sinef <= -565;
 when 2094 => sinef <= -578;
 when 2095 => sinef <= -590;
 when 2096 => sinef <= -603;
 when 2097 => sinef <= -615;
 when 2098 => sinef <= -628;
 when 2099 => sinef <= -640;
 when 2100 => sinef <= -653;
 when 2101 => sinef <= -665;
 when 2102 => sinef <= -678;
 when 2103 => sinef <= -690;
 when 2104 => sinef <= -703;
 when 2105 => sinef <= -715;
 when 2106 => sinef <= -728;
 when 2107 => sinef <= -740;
 when 2108 => sinef <= -753;
 when 2109 => sinef <= -765;
 when 2110 => sinef <= -778;
 when 2111 => sinef <= -790;
 when 2112 => sinef <= -803;
 when 2113 => sinef <= -815;
 when 2114 => sinef <= -828;
 when 2115 => sinef <= -840;
 when 2116 => sinef <= -853;
 when 2117 => sinef <= -865;
 when 2118 => sinef <= -878;
 when 2119 => sinef <= -890;
 when 2120 => sinef <= -903;
 when 2121 => sinef <= -915;
 when 2122 => sinef <= -928;
 when 2123 => sinef <= -940;
 when 2124 => sinef <= -953;
 when 2125 => sinef <= -965;
 when 2126 => sinef <= -978;
 when 2127 => sinef <= -990;
 when 2128 => sinef <= -1003;
 when 2129 => sinef <= -1015;
 when 2130 => sinef <= -1028;
 when 2131 => sinef <= -1040;
 when 2132 => sinef <= -1053;
 when 2133 => sinef <= -1065;
 when 2134 => sinef <= -1077;
 when 2135 => sinef <= -1090;
 when 2136 => sinef <= -1102;
 when 2137 => sinef <= -1115;
 when 2138 => sinef <= -1127;
 when 2139 => sinef <= -1140;
 when 2140 => sinef <= -1152;
 when 2141 => sinef <= -1165;
 when 2142 => sinef <= -1177;
 when 2143 => sinef <= -1189;
 when 2144 => sinef <= -1202;
 when 2145 => sinef <= -1214;
 when 2146 => sinef <= -1227;
 when 2147 => sinef <= -1239;
 when 2148 => sinef <= -1252;
 when 2149 => sinef <= -1264;
 when 2150 => sinef <= -1276;
 when 2151 => sinef <= -1289;
 when 2152 => sinef <= -1301;
 when 2153 => sinef <= -1314;
 when 2154 => sinef <= -1326;
 when 2155 => sinef <= -1338;
 when 2156 => sinef <= -1351;
 when 2157 => sinef <= -1363;
 when 2158 => sinef <= -1376;
 when 2159 => sinef <= -1388;
 when 2160 => sinef <= -1400;
 when 2161 => sinef <= -1413;
 when 2162 => sinef <= -1425;
 when 2163 => sinef <= -1437;
 when 2164 => sinef <= -1450;
 when 2165 => sinef <= -1462;
 when 2166 => sinef <= -1475;
 when 2167 => sinef <= -1487;
 when 2168 => sinef <= -1499;
 when 2169 => sinef <= -1512;
 when 2170 => sinef <= -1524;
 when 2171 => sinef <= -1536;
 when 2172 => sinef <= -1549;
 when 2173 => sinef <= -1561;
 when 2174 => sinef <= -1573;
 when 2175 => sinef <= -1586;
 when 2176 => sinef <= -1598;
 when 2177 => sinef <= -1610;
 when 2178 => sinef <= -1623;
 when 2179 => sinef <= -1635;
 when 2180 => sinef <= -1647;
 when 2181 => sinef <= -1660;
 when 2182 => sinef <= -1672;
 when 2183 => sinef <= -1684;
 when 2184 => sinef <= -1696;
 when 2185 => sinef <= -1709;
 when 2186 => sinef <= -1721;
 when 2187 => sinef <= -1733;
 when 2188 => sinef <= -1746;
 when 2189 => sinef <= -1758;
 when 2190 => sinef <= -1770;
 when 2191 => sinef <= -1782;
 when 2192 => sinef <= -1795;
 when 2193 => sinef <= -1807;
 when 2194 => sinef <= -1819;
 when 2195 => sinef <= -1831;
 when 2196 => sinef <= -1844;
 when 2197 => sinef <= -1856;
 when 2198 => sinef <= -1868;
 when 2199 => sinef <= -1880;
 when 2200 => sinef <= -1893;
 when 2201 => sinef <= -1905;
 when 2202 => sinef <= -1917;
 when 2203 => sinef <= -1929;
 when 2204 => sinef <= -1941;
 when 2205 => sinef <= -1954;
 when 2206 => sinef <= -1966;
 when 2207 => sinef <= -1978;
 when 2208 => sinef <= -1990;
 when 2209 => sinef <= -2002;
 when 2210 => sinef <= -2015;
 when 2211 => sinef <= -2027;
 when 2212 => sinef <= -2039;
 when 2213 => sinef <= -2051;
 when 2214 => sinef <= -2063;
 when 2215 => sinef <= -2075;
 when 2216 => sinef <= -2088;
 when 2217 => sinef <= -2100;
 when 2218 => sinef <= -2112;
 when 2219 => sinef <= -2124;
 when 2220 => sinef <= -2136;
 when 2221 => sinef <= -2148;
 when 2222 => sinef <= -2160;
 when 2223 => sinef <= -2173;
 when 2224 => sinef <= -2185;
 when 2225 => sinef <= -2197;
 when 2226 => sinef <= -2209;
 when 2227 => sinef <= -2221;
 when 2228 => sinef <= -2233;
 when 2229 => sinef <= -2245;
 when 2230 => sinef <= -2257;
 when 2231 => sinef <= -2269;
 when 2232 => sinef <= -2281;
 when 2233 => sinef <= -2293;
 when 2234 => sinef <= -2305;
 when 2235 => sinef <= -2318;
 when 2236 => sinef <= -2330;
 when 2237 => sinef <= -2342;
 when 2238 => sinef <= -2354;
 when 2239 => sinef <= -2366;
 when 2240 => sinef <= -2378;
 when 2241 => sinef <= -2390;
 when 2242 => sinef <= -2402;
 when 2243 => sinef <= -2414;
 when 2244 => sinef <= -2426;
 when 2245 => sinef <= -2438;
 when 2246 => sinef <= -2450;
 when 2247 => sinef <= -2462;
 when 2248 => sinef <= -2474;
 when 2249 => sinef <= -2486;
 when 2250 => sinef <= -2498;
 when 2251 => sinef <= -2510;
 when 2252 => sinef <= -2522;
 when 2253 => sinef <= -2534;
 when 2254 => sinef <= -2545;
 when 2255 => sinef <= -2557;
 when 2256 => sinef <= -2569;
 when 2257 => sinef <= -2581;
 when 2258 => sinef <= -2593;
 when 2259 => sinef <= -2605;
 when 2260 => sinef <= -2617;
 when 2261 => sinef <= -2629;
 when 2262 => sinef <= -2641;
 when 2263 => sinef <= -2653;
 when 2264 => sinef <= -2665;
 when 2265 => sinef <= -2676;
 when 2266 => sinef <= -2688;
 when 2267 => sinef <= -2700;
 when 2268 => sinef <= -2712;
 when 2269 => sinef <= -2724;
 when 2270 => sinef <= -2736;
 when 2271 => sinef <= -2748;
 when 2272 => sinef <= -2759;
 when 2273 => sinef <= -2771;
 when 2274 => sinef <= -2783;
 when 2275 => sinef <= -2795;
 when 2276 => sinef <= -2807;
 when 2277 => sinef <= -2819;
 when 2278 => sinef <= -2830;
 when 2279 => sinef <= -2842;
 when 2280 => sinef <= -2854;
 when 2281 => sinef <= -2866;
 when 2282 => sinef <= -2877;
 when 2283 => sinef <= -2889;
 when 2284 => sinef <= -2901;
 when 2285 => sinef <= -2913;
 when 2286 => sinef <= -2924;
 when 2287 => sinef <= -2936;
 when 2288 => sinef <= -2948;
 when 2289 => sinef <= -2960;
 when 2290 => sinef <= -2971;
 when 2291 => sinef <= -2983;
 when 2292 => sinef <= -2995;
 when 2293 => sinef <= -3006;
 when 2294 => sinef <= -3018;
 when 2295 => sinef <= -3030;
 when 2296 => sinef <= -3041;
 when 2297 => sinef <= -3053;
 when 2298 => sinef <= -3065;
 when 2299 => sinef <= -3076;
 when 2300 => sinef <= -3088;
 when 2301 => sinef <= -3100;
 when 2302 => sinef <= -3111;
 when 2303 => sinef <= -3123;
 when 2304 => sinef <= -3135;
 when 2305 => sinef <= -3146;
 when 2306 => sinef <= -3158;
 when 2307 => sinef <= -3169;
 when 2308 => sinef <= -3181;
 when 2309 => sinef <= -3193;
 when 2310 => sinef <= -3204;
 when 2311 => sinef <= -3216;
 when 2312 => sinef <= -3227;
 when 2313 => sinef <= -3239;
 when 2314 => sinef <= -3250;
 when 2315 => sinef <= -3262;
 when 2316 => sinef <= -3273;
 when 2317 => sinef <= -3285;
 when 2318 => sinef <= -3296;
 when 2319 => sinef <= -3308;
 when 2320 => sinef <= -3319;
 when 2321 => sinef <= -3331;
 when 2322 => sinef <= -3342;
 when 2323 => sinef <= -3354;
 when 2324 => sinef <= -3365;
 when 2325 => sinef <= -3377;
 when 2326 => sinef <= -3388;
 when 2327 => sinef <= -3400;
 when 2328 => sinef <= -3411;
 when 2329 => sinef <= -3422;
 when 2330 => sinef <= -3434;
 when 2331 => sinef <= -3445;
 when 2332 => sinef <= -3457;
 when 2333 => sinef <= -3468;
 when 2334 => sinef <= -3479;
 when 2335 => sinef <= -3491;
 when 2336 => sinef <= -3502;
 when 2337 => sinef <= -3513;
 when 2338 => sinef <= -3525;
 when 2339 => sinef <= -3536;
 when 2340 => sinef <= -3547;
 when 2341 => sinef <= -3559;
 when 2342 => sinef <= -3570;
 when 2343 => sinef <= -3581;
 when 2344 => sinef <= -3593;
 when 2345 => sinef <= -3604;
 when 2346 => sinef <= -3615;
 when 2347 => sinef <= -3627;
 when 2348 => sinef <= -3638;
 when 2349 => sinef <= -3649;
 when 2350 => sinef <= -3660;
 when 2351 => sinef <= -3672;
 when 2352 => sinef <= -3683;
 when 2353 => sinef <= -3694;
 when 2354 => sinef <= -3705;
 when 2355 => sinef <= -3716;
 when 2356 => sinef <= -3728;
 when 2357 => sinef <= -3739;
 when 2358 => sinef <= -3750;
 when 2359 => sinef <= -3761;
 when 2360 => sinef <= -3772;
 when 2361 => sinef <= -3783;
 when 2362 => sinef <= -3795;
 when 2363 => sinef <= -3806;
 when 2364 => sinef <= -3817;
 when 2365 => sinef <= -3828;
 when 2366 => sinef <= -3839;
 when 2367 => sinef <= -3850;
 when 2368 => sinef <= -3861;
 when 2369 => sinef <= -3872;
 when 2370 => sinef <= -3883;
 when 2371 => sinef <= -3894;
 when 2372 => sinef <= -3905;
 when 2373 => sinef <= -3917;
 when 2374 => sinef <= -3928;
 when 2375 => sinef <= -3939;
 when 2376 => sinef <= -3950;
 when 2377 => sinef <= -3961;
 when 2378 => sinef <= -3972;
 when 2379 => sinef <= -3983;
 when 2380 => sinef <= -3994;
 when 2381 => sinef <= -4004;
 when 2382 => sinef <= -4015;
 when 2383 => sinef <= -4026;
 when 2384 => sinef <= -4037;
 when 2385 => sinef <= -4048;
 when 2386 => sinef <= -4059;
 when 2387 => sinef <= -4070;
 when 2388 => sinef <= -4081;
 when 2389 => sinef <= -4092;
 when 2390 => sinef <= -4103;
 when 2391 => sinef <= -4114;
 when 2392 => sinef <= -4124;
 when 2393 => sinef <= -4135;
 when 2394 => sinef <= -4146;
 when 2395 => sinef <= -4157;
 when 2396 => sinef <= -4168;
 when 2397 => sinef <= -4179;
 when 2398 => sinef <= -4189;
 when 2399 => sinef <= -4200;
 when 2400 => sinef <= -4211;
 when 2401 => sinef <= -4222;
 when 2402 => sinef <= -4233;
 when 2403 => sinef <= -4243;
 when 2404 => sinef <= -4254;
 when 2405 => sinef <= -4265;
 when 2406 => sinef <= -4275;
 when 2407 => sinef <= -4286;
 when 2408 => sinef <= -4297;
 when 2409 => sinef <= -4308;
 when 2410 => sinef <= -4318;
 when 2411 => sinef <= -4329;
 when 2412 => sinef <= -4340;
 when 2413 => sinef <= -4350;
 when 2414 => sinef <= -4361;
 when 2415 => sinef <= -4372;
 when 2416 => sinef <= -4382;
 when 2417 => sinef <= -4393;
 when 2418 => sinef <= -4403;
 when 2419 => sinef <= -4414;
 when 2420 => sinef <= -4425;
 when 2421 => sinef <= -4435;
 when 2422 => sinef <= -4446;
 when 2423 => sinef <= -4456;
 when 2424 => sinef <= -4467;
 when 2425 => sinef <= -4477;
 when 2426 => sinef <= -4488;
 when 2427 => sinef <= -4498;
 when 2428 => sinef <= -4509;
 when 2429 => sinef <= -4519;
 when 2430 => sinef <= -4530;
 when 2431 => sinef <= -4540;
 when 2432 => sinef <= -4551;
 when 2433 => sinef <= -4561;
 when 2434 => sinef <= -4572;
 when 2435 => sinef <= -4582;
 when 2436 => sinef <= -4592;
 when 2437 => sinef <= -4603;
 when 2438 => sinef <= -4613;
 when 2439 => sinef <= -4624;
 when 2440 => sinef <= -4634;
 when 2441 => sinef <= -4644;
 when 2442 => sinef <= -4655;
 when 2443 => sinef <= -4665;
 when 2444 => sinef <= -4675;
 when 2445 => sinef <= -4686;
 when 2446 => sinef <= -4696;
 when 2447 => sinef <= -4706;
 when 2448 => sinef <= -4716;
 when 2449 => sinef <= -4727;
 when 2450 => sinef <= -4737;
 when 2451 => sinef <= -4747;
 when 2452 => sinef <= -4757;
 when 2453 => sinef <= -4768;
 when 2454 => sinef <= -4778;
 when 2455 => sinef <= -4788;
 when 2456 => sinef <= -4798;
 when 2457 => sinef <= -4808;
 when 2458 => sinef <= -4819;
 when 2459 => sinef <= -4829;
 when 2460 => sinef <= -4839;
 when 2461 => sinef <= -4849;
 when 2462 => sinef <= -4859;
 when 2463 => sinef <= -4869;
 when 2464 => sinef <= -4879;
 when 2465 => sinef <= -4889;
 when 2466 => sinef <= -4900;
 when 2467 => sinef <= -4910;
 when 2468 => sinef <= -4920;
 when 2469 => sinef <= -4930;
 when 2470 => sinef <= -4940;
 when 2471 => sinef <= -4950;
 when 2472 => sinef <= -4960;
 when 2473 => sinef <= -4970;
 when 2474 => sinef <= -4980;
 when 2475 => sinef <= -4990;
 when 2476 => sinef <= -5000;
 when 2477 => sinef <= -5010;
 when 2478 => sinef <= -5020;
 when 2479 => sinef <= -5029;
 when 2480 => sinef <= -5039;
 when 2481 => sinef <= -5049;
 when 2482 => sinef <= -5059;
 when 2483 => sinef <= -5069;
 when 2484 => sinef <= -5079;
 when 2485 => sinef <= -5089;
 when 2486 => sinef <= -5099;
 when 2487 => sinef <= -5108;
 when 2488 => sinef <= -5118;
 when 2489 => sinef <= -5128;
 when 2490 => sinef <= -5138;
 when 2491 => sinef <= -5148;
 when 2492 => sinef <= -5157;
 when 2493 => sinef <= -5167;
 when 2494 => sinef <= -5177;
 when 2495 => sinef <= -5187;
 when 2496 => sinef <= -5196;
 when 2497 => sinef <= -5206;
 when 2498 => sinef <= -5216;
 when 2499 => sinef <= -5225;
 when 2500 => sinef <= -5235;
 when 2501 => sinef <= -5245;
 when 2502 => sinef <= -5254;
 when 2503 => sinef <= -5264;
 when 2504 => sinef <= -5274;
 when 2505 => sinef <= -5283;
 when 2506 => sinef <= -5293;
 when 2507 => sinef <= -5302;
 when 2508 => sinef <= -5312;
 when 2509 => sinef <= -5322;
 when 2510 => sinef <= -5331;
 when 2511 => sinef <= -5341;
 when 2512 => sinef <= -5350;
 when 2513 => sinef <= -5360;
 when 2514 => sinef <= -5369;
 when 2515 => sinef <= -5379;
 when 2516 => sinef <= -5388;
 when 2517 => sinef <= -5398;
 when 2518 => sinef <= -5407;
 when 2519 => sinef <= -5416;
 when 2520 => sinef <= -5426;
 when 2521 => sinef <= -5435;
 when 2522 => sinef <= -5445;
 when 2523 => sinef <= -5454;
 when 2524 => sinef <= -5463;
 when 2525 => sinef <= -5473;
 when 2526 => sinef <= -5482;
 when 2527 => sinef <= -5491;
 when 2528 => sinef <= -5501;
 when 2529 => sinef <= -5510;
 when 2530 => sinef <= -5519;
 when 2531 => sinef <= -5529;
 when 2532 => sinef <= -5538;
 when 2533 => sinef <= -5547;
 when 2534 => sinef <= -5556;
 when 2535 => sinef <= -5566;
 when 2536 => sinef <= -5575;
 when 2537 => sinef <= -5584;
 when 2538 => sinef <= -5593;
 when 2539 => sinef <= -5602;
 when 2540 => sinef <= -5612;
 when 2541 => sinef <= -5621;
 when 2542 => sinef <= -5630;
 when 2543 => sinef <= -5639;
 when 2544 => sinef <= -5648;
 when 2545 => sinef <= -5657;
 when 2546 => sinef <= -5666;
 when 2547 => sinef <= -5675;
 when 2548 => sinef <= -5684;
 when 2549 => sinef <= -5693;
 when 2550 => sinef <= -5702;
 when 2551 => sinef <= -5711;
 when 2552 => sinef <= -5720;
 when 2553 => sinef <= -5729;
 when 2554 => sinef <= -5738;
 when 2555 => sinef <= -5747;
 when 2556 => sinef <= -5756;
 when 2557 => sinef <= -5765;
 when 2558 => sinef <= -5774;
 when 2559 => sinef <= -5783;
 when 2560 => sinef <= -5792;
 when 2561 => sinef <= -5801;
 when 2562 => sinef <= -5810;
 when 2563 => sinef <= -5819;
 when 2564 => sinef <= -5827;
 when 2565 => sinef <= -5836;
 when 2566 => sinef <= -5845;
 when 2567 => sinef <= -5854;
 when 2568 => sinef <= -5863;
 when 2569 => sinef <= -5871;
 when 2570 => sinef <= -5880;
 when 2571 => sinef <= -5889;
 when 2572 => sinef <= -5898;
 when 2573 => sinef <= -5906;
 when 2574 => sinef <= -5915;
 when 2575 => sinef <= -5924;
 when 2576 => sinef <= -5932;
 when 2577 => sinef <= -5941;
 when 2578 => sinef <= -5950;
 when 2579 => sinef <= -5958;
 when 2580 => sinef <= -5967;
 when 2581 => sinef <= -5975;
 when 2582 => sinef <= -5984;
 when 2583 => sinef <= -5993;
 when 2584 => sinef <= -6001;
 when 2585 => sinef <= -6010;
 when 2586 => sinef <= -6018;
 when 2587 => sinef <= -6027;
 when 2588 => sinef <= -6035;
 when 2589 => sinef <= -6044;
 when 2590 => sinef <= -6052;
 when 2591 => sinef <= -6061;
 when 2592 => sinef <= -6069;
 when 2593 => sinef <= -6078;
 when 2594 => sinef <= -6086;
 when 2595 => sinef <= -6094;
 when 2596 => sinef <= -6103;
 when 2597 => sinef <= -6111;
 when 2598 => sinef <= -6120;
 when 2599 => sinef <= -6128;
 when 2600 => sinef <= -6136;
 when 2601 => sinef <= -6144;
 when 2602 => sinef <= -6153;
 when 2603 => sinef <= -6161;
 when 2604 => sinef <= -6169;
 when 2605 => sinef <= -6178;
 when 2606 => sinef <= -6186;
 when 2607 => sinef <= -6194;
 when 2608 => sinef <= -6202;
 when 2609 => sinef <= -6210;
 when 2610 => sinef <= -6219;
 when 2611 => sinef <= -6227;
 when 2612 => sinef <= -6235;
 when 2613 => sinef <= -6243;
 when 2614 => sinef <= -6251;
 when 2615 => sinef <= -6259;
 when 2616 => sinef <= -6267;
 when 2617 => sinef <= -6276;
 when 2618 => sinef <= -6284;
 when 2619 => sinef <= -6292;
 when 2620 => sinef <= -6300;
 when 2621 => sinef <= -6308;
 when 2622 => sinef <= -6316;
 when 2623 => sinef <= -6324;
 when 2624 => sinef <= -6332;
 when 2625 => sinef <= -6340;
 when 2626 => sinef <= -6348;
 when 2627 => sinef <= -6356;
 when 2628 => sinef <= -6363;
 when 2629 => sinef <= -6371;
 when 2630 => sinef <= -6379;
 when 2631 => sinef <= -6387;
 when 2632 => sinef <= -6395;
 when 2633 => sinef <= -6403;
 when 2634 => sinef <= -6411;
 when 2635 => sinef <= -6419;
 when 2636 => sinef <= -6426;
 when 2637 => sinef <= -6434;
 when 2638 => sinef <= -6442;
 when 2639 => sinef <= -6450;
 when 2640 => sinef <= -6457;
 when 2641 => sinef <= -6465;
 when 2642 => sinef <= -6473;
 when 2643 => sinef <= -6480;
 when 2644 => sinef <= -6488;
 when 2645 => sinef <= -6496;
 when 2646 => sinef <= -6503;
 when 2647 => sinef <= -6511;
 when 2648 => sinef <= -6519;
 when 2649 => sinef <= -6526;
 when 2650 => sinef <= -6534;
 when 2651 => sinef <= -6541;
 when 2652 => sinef <= -6549;
 when 2653 => sinef <= -6557;
 when 2654 => sinef <= -6564;
 when 2655 => sinef <= -6572;
 when 2656 => sinef <= -6579;
 when 2657 => sinef <= -6587;
 when 2658 => sinef <= -6594;
 when 2659 => sinef <= -6601;
 when 2660 => sinef <= -6609;
 when 2661 => sinef <= -6616;
 when 2662 => sinef <= -6624;
 when 2663 => sinef <= -6631;
 when 2664 => sinef <= -6638;
 when 2665 => sinef <= -6646;
 when 2666 => sinef <= -6653;
 when 2667 => sinef <= -6660;
 when 2668 => sinef <= -6668;
 when 2669 => sinef <= -6675;
 when 2670 => sinef <= -6682;
 when 2671 => sinef <= -6690;
 when 2672 => sinef <= -6697;
 when 2673 => sinef <= -6704;
 when 2674 => sinef <= -6711;
 when 2675 => sinef <= -6718;
 when 2676 => sinef <= -6726;
 when 2677 => sinef <= -6733;
 when 2678 => sinef <= -6740;
 when 2679 => sinef <= -6747;
 when 2680 => sinef <= -6754;
 when 2681 => sinef <= -6761;
 when 2682 => sinef <= -6768;
 when 2683 => sinef <= -6775;
 when 2684 => sinef <= -6783;
 when 2685 => sinef <= -6790;
 when 2686 => sinef <= -6797;
 when 2687 => sinef <= -6804;
 when 2688 => sinef <= -6811;
 when 2689 => sinef <= -6818;
 when 2690 => sinef <= -6824;
 when 2691 => sinef <= -6831;
 when 2692 => sinef <= -6838;
 when 2693 => sinef <= -6845;
 when 2694 => sinef <= -6852;
 when 2695 => sinef <= -6859;
 when 2696 => sinef <= -6866;
 when 2697 => sinef <= -6873;
 when 2698 => sinef <= -6880;
 when 2699 => sinef <= -6886;
 when 2700 => sinef <= -6893;
 when 2701 => sinef <= -6900;
 when 2702 => sinef <= -6907;
 when 2703 => sinef <= -6913;
 when 2704 => sinef <= -6920;
 when 2705 => sinef <= -6927;
 when 2706 => sinef <= -6934;
 when 2707 => sinef <= -6940;
 when 2708 => sinef <= -6947;
 when 2709 => sinef <= -6954;
 when 2710 => sinef <= -6960;
 when 2711 => sinef <= -6967;
 when 2712 => sinef <= -6973;
 when 2713 => sinef <= -6980;
 when 2714 => sinef <= -6987;
 when 2715 => sinef <= -6993;
 when 2716 => sinef <= -7000;
 when 2717 => sinef <= -7006;
 when 2718 => sinef <= -7013;
 when 2719 => sinef <= -7019;
 when 2720 => sinef <= -7026;
 when 2721 => sinef <= -7032;
 when 2722 => sinef <= -7039;
 when 2723 => sinef <= -7045;
 when 2724 => sinef <= -7051;
 when 2725 => sinef <= -7058;
 when 2726 => sinef <= -7064;
 when 2727 => sinef <= -7070;
 when 2728 => sinef <= -7077;
 when 2729 => sinef <= -7083;
 when 2730 => sinef <= -7089;
 when 2731 => sinef <= -7096;
 when 2732 => sinef <= -7102;
 when 2733 => sinef <= -7108;
 when 2734 => sinef <= -7114;
 when 2735 => sinef <= -7121;
 when 2736 => sinef <= -7127;
 when 2737 => sinef <= -7133;
 when 2738 => sinef <= -7139;
 when 2739 => sinef <= -7145;
 when 2740 => sinef <= -7152;
 when 2741 => sinef <= -7158;
 when 2742 => sinef <= -7164;
 when 2743 => sinef <= -7170;
 when 2744 => sinef <= -7176;
 when 2745 => sinef <= -7182;
 when 2746 => sinef <= -7188;
 when 2747 => sinef <= -7194;
 when 2748 => sinef <= -7200;
 when 2749 => sinef <= -7206;
 when 2750 => sinef <= -7212;
 when 2751 => sinef <= -7218;
 when 2752 => sinef <= -7224;
 when 2753 => sinef <= -7230;
 when 2754 => sinef <= -7236;
 when 2755 => sinef <= -7242;
 when 2756 => sinef <= -7247;
 when 2757 => sinef <= -7253;
 when 2758 => sinef <= -7259;
 when 2759 => sinef <= -7265;
 when 2760 => sinef <= -7271;
 when 2761 => sinef <= -7276;
 when 2762 => sinef <= -7282;
 when 2763 => sinef <= -7288;
 when 2764 => sinef <= -7294;
 when 2765 => sinef <= -7299;
 when 2766 => sinef <= -7305;
 when 2767 => sinef <= -7311;
 when 2768 => sinef <= -7316;
 when 2769 => sinef <= -7322;
 when 2770 => sinef <= -7328;
 when 2771 => sinef <= -7333;
 when 2772 => sinef <= -7339;
 when 2773 => sinef <= -7344;
 when 2774 => sinef <= -7350;
 when 2775 => sinef <= -7356;
 when 2776 => sinef <= -7361;
 when 2777 => sinef <= -7367;
 when 2778 => sinef <= -7372;
 when 2779 => sinef <= -7377;
 when 2780 => sinef <= -7383;
 when 2781 => sinef <= -7388;
 when 2782 => sinef <= -7394;
 when 2783 => sinef <= -7399;
 when 2784 => sinef <= -7405;
 when 2785 => sinef <= -7410;
 when 2786 => sinef <= -7415;
 when 2787 => sinef <= -7421;
 when 2788 => sinef <= -7426;
 when 2789 => sinef <= -7431;
 when 2790 => sinef <= -7436;
 when 2791 => sinef <= -7442;
 when 2792 => sinef <= -7447;
 when 2793 => sinef <= -7452;
 when 2794 => sinef <= -7457;
 when 2795 => sinef <= -7463;
 when 2796 => sinef <= -7468;
 when 2797 => sinef <= -7473;
 when 2798 => sinef <= -7478;
 when 2799 => sinef <= -7483;
 when 2800 => sinef <= -7488;
 when 2801 => sinef <= -7493;
 when 2802 => sinef <= -7498;
 when 2803 => sinef <= -7503;
 when 2804 => sinef <= -7509;
 when 2805 => sinef <= -7514;
 when 2806 => sinef <= -7519;
 when 2807 => sinef <= -7524;
 when 2808 => sinef <= -7528;
 when 2809 => sinef <= -7533;
 when 2810 => sinef <= -7538;
 when 2811 => sinef <= -7543;
 when 2812 => sinef <= -7548;
 when 2813 => sinef <= -7553;
 when 2814 => sinef <= -7558;
 when 2815 => sinef <= -7563;
 when 2816 => sinef <= -7567;
 when 2817 => sinef <= -7572;
 when 2818 => sinef <= -7577;
 when 2819 => sinef <= -7582;
 when 2820 => sinef <= -7587;
 when 2821 => sinef <= -7591;
 when 2822 => sinef <= -7596;
 when 2823 => sinef <= -7601;
 when 2824 => sinef <= -7605;
 when 2825 => sinef <= -7610;
 when 2826 => sinef <= -7615;
 when 2827 => sinef <= -7619;
 when 2828 => sinef <= -7624;
 when 2829 => sinef <= -7628;
 when 2830 => sinef <= -7633;
 when 2831 => sinef <= -7638;
 when 2832 => sinef <= -7642;
 when 2833 => sinef <= -7647;
 when 2834 => sinef <= -7651;
 when 2835 => sinef <= -7656;
 when 2836 => sinef <= -7660;
 when 2837 => sinef <= -7665;
 when 2838 => sinef <= -7669;
 when 2839 => sinef <= -7673;
 when 2840 => sinef <= -7678;
 when 2841 => sinef <= -7682;
 when 2842 => sinef <= -7686;
 when 2843 => sinef <= -7691;
 when 2844 => sinef <= -7695;
 when 2845 => sinef <= -7699;
 when 2846 => sinef <= -7704;
 when 2847 => sinef <= -7708;
 when 2848 => sinef <= -7712;
 when 2849 => sinef <= -7716;
 when 2850 => sinef <= -7721;
 when 2851 => sinef <= -7725;
 when 2852 => sinef <= -7729;
 when 2853 => sinef <= -7733;
 when 2854 => sinef <= -7737;
 when 2855 => sinef <= -7741;
 when 2856 => sinef <= -7745;
 when 2857 => sinef <= -7750;
 when 2858 => sinef <= -7754;
 when 2859 => sinef <= -7758;
 when 2860 => sinef <= -7762;
 when 2861 => sinef <= -7766;
 when 2862 => sinef <= -7770;
 when 2863 => sinef <= -7774;
 when 2864 => sinef <= -7778;
 when 2865 => sinef <= -7782;
 when 2866 => sinef <= -7785;
 when 2867 => sinef <= -7789;
 when 2868 => sinef <= -7793;
 when 2869 => sinef <= -7797;
 when 2870 => sinef <= -7801;
 when 2871 => sinef <= -7805;
 when 2872 => sinef <= -7809;
 when 2873 => sinef <= -7812;
 when 2874 => sinef <= -7816;
 when 2875 => sinef <= -7820;
 when 2876 => sinef <= -7824;
 when 2877 => sinef <= -7827;
 when 2878 => sinef <= -7831;
 when 2879 => sinef <= -7835;
 when 2880 => sinef <= -7838;
 when 2881 => sinef <= -7842;
 when 2882 => sinef <= -7846;
 when 2883 => sinef <= -7849;
 when 2884 => sinef <= -7853;
 when 2885 => sinef <= -7856;
 when 2886 => sinef <= -7860;
 when 2887 => sinef <= -7863;
 when 2888 => sinef <= -7867;
 when 2889 => sinef <= -7870;
 when 2890 => sinef <= -7874;
 when 2891 => sinef <= -7877;
 when 2892 => sinef <= -7881;
 when 2893 => sinef <= -7884;
 when 2894 => sinef <= -7888;
 when 2895 => sinef <= -7891;
 when 2896 => sinef <= -7894;
 when 2897 => sinef <= -7898;
 when 2898 => sinef <= -7901;
 when 2899 => sinef <= -7904;
 when 2900 => sinef <= -7908;
 when 2901 => sinef <= -7911;
 when 2902 => sinef <= -7914;
 when 2903 => sinef <= -7917;
 when 2904 => sinef <= -7921;
 when 2905 => sinef <= -7924;
 when 2906 => sinef <= -7927;
 when 2907 => sinef <= -7930;
 when 2908 => sinef <= -7933;
 when 2909 => sinef <= -7936;
 when 2910 => sinef <= -7939;
 when 2911 => sinef <= -7942;
 when 2912 => sinef <= -7946;
 when 2913 => sinef <= -7949;
 when 2914 => sinef <= -7952;
 when 2915 => sinef <= -7955;
 when 2916 => sinef <= -7958;
 when 2917 => sinef <= -7961;
 when 2918 => sinef <= -7964;
 when 2919 => sinef <= -7966;
 when 2920 => sinef <= -7969;
 when 2921 => sinef <= -7972;
 when 2922 => sinef <= -7975;
 when 2923 => sinef <= -7978;
 when 2924 => sinef <= -7981;
 when 2925 => sinef <= -7984;
 when 2926 => sinef <= -7986;
 when 2927 => sinef <= -7989;
 when 2928 => sinef <= -7992;
 when 2929 => sinef <= -7995;
 when 2930 => sinef <= -7997;
 when 2931 => sinef <= -8000;
 when 2932 => sinef <= -8003;
 when 2933 => sinef <= -8006;
 when 2934 => sinef <= -8008;
 when 2935 => sinef <= -8011;
 when 2936 => sinef <= -8013;
 when 2937 => sinef <= -8016;
 when 2938 => sinef <= -8019;
 when 2939 => sinef <= -8021;
 when 2940 => sinef <= -8024;
 when 2941 => sinef <= -8026;
 when 2942 => sinef <= -8029;
 when 2943 => sinef <= -8031;
 when 2944 => sinef <= -8034;
 when 2945 => sinef <= -8036;
 when 2946 => sinef <= -8038;
 when 2947 => sinef <= -8041;
 when 2948 => sinef <= -8043;
 when 2949 => sinef <= -8046;
 when 2950 => sinef <= -8048;
 when 2951 => sinef <= -8050;
 when 2952 => sinef <= -8053;
 when 2953 => sinef <= -8055;
 when 2954 => sinef <= -8057;
 when 2955 => sinef <= -8059;
 when 2956 => sinef <= -8062;
 when 2957 => sinef <= -8064;
 when 2958 => sinef <= -8066;
 when 2959 => sinef <= -8068;
 when 2960 => sinef <= -8070;
 when 2961 => sinef <= -8073;
 when 2962 => sinef <= -8075;
 when 2963 => sinef <= -8077;
 when 2964 => sinef <= -8079;
 when 2965 => sinef <= -8081;
 when 2966 => sinef <= -8083;
 when 2967 => sinef <= -8085;
 when 2968 => sinef <= -8087;
 when 2969 => sinef <= -8089;
 when 2970 => sinef <= -8091;
 when 2971 => sinef <= -8093;
 when 2972 => sinef <= -8095;
 when 2973 => sinef <= -8097;
 when 2974 => sinef <= -8099;
 when 2975 => sinef <= -8100;
 when 2976 => sinef <= -8102;
 when 2977 => sinef <= -8104;
 when 2978 => sinef <= -8106;
 when 2979 => sinef <= -8108;
 when 2980 => sinef <= -8110;
 when 2981 => sinef <= -8111;
 when 2982 => sinef <= -8113;
 when 2983 => sinef <= -8115;
 when 2984 => sinef <= -8116;
 when 2985 => sinef <= -8118;
 when 2986 => sinef <= -8120;
 when 2987 => sinef <= -8121;
 when 2988 => sinef <= -8123;
 when 2989 => sinef <= -8125;
 when 2990 => sinef <= -8126;
 when 2991 => sinef <= -8128;
 when 2992 => sinef <= -8129;
 when 2993 => sinef <= -8131;
 when 2994 => sinef <= -8132;
 when 2995 => sinef <= -8134;
 when 2996 => sinef <= -8135;
 when 2997 => sinef <= -8137;
 when 2998 => sinef <= -8138;
 when 2999 => sinef <= -8140;
 when 3000 => sinef <= -8141;
 when 3001 => sinef <= -8142;
 when 3002 => sinef <= -8144;
 when 3003 => sinef <= -8145;
 when 3004 => sinef <= -8146;
 when 3005 => sinef <= -8148;
 when 3006 => sinef <= -8149;
 when 3007 => sinef <= -8150;
 when 3008 => sinef <= -8152;
 when 3009 => sinef <= -8153;
 when 3010 => sinef <= -8154;
 when 3011 => sinef <= -8155;
 when 3012 => sinef <= -8156;
 when 3013 => sinef <= -8157;
 when 3014 => sinef <= -8159;
 when 3015 => sinef <= -8160;
 when 3016 => sinef <= -8161;
 when 3017 => sinef <= -8162;
 when 3018 => sinef <= -8163;
 when 3019 => sinef <= -8164;
 when 3020 => sinef <= -8165;
 when 3021 => sinef <= -8166;
 when 3022 => sinef <= -8167;
 when 3023 => sinef <= -8168;
 when 3024 => sinef <= -8169;
 when 3025 => sinef <= -8170;
 when 3026 => sinef <= -8171;
 when 3027 => sinef <= -8171;
 when 3028 => sinef <= -8172;
 when 3029 => sinef <= -8173;
 when 3030 => sinef <= -8174;
 when 3031 => sinef <= -8175;
 when 3032 => sinef <= -8176;
 when 3033 => sinef <= -8176;
 when 3034 => sinef <= -8177;
 when 3035 => sinef <= -8178;
 when 3036 => sinef <= -8179;
 when 3037 => sinef <= -8179;
 when 3038 => sinef <= -8180;
 when 3039 => sinef <= -8181;
 when 3040 => sinef <= -8181;
 when 3041 => sinef <= -8182;
 when 3042 => sinef <= -8182;
 when 3043 => sinef <= -8183;
 when 3044 => sinef <= -8183;
 when 3045 => sinef <= -8184;
 when 3046 => sinef <= -8184;
 when 3047 => sinef <= -8185;
 when 3048 => sinef <= -8185;
 when 3049 => sinef <= -8186;
 when 3050 => sinef <= -8186;
 when 3051 => sinef <= -8187;
 when 3052 => sinef <= -8187;
 when 3053 => sinef <= -8188;
 when 3054 => sinef <= -8188;
 when 3055 => sinef <= -8188;
 when 3056 => sinef <= -8189;
 when 3057 => sinef <= -8189;
 when 3058 => sinef <= -8189;
 when 3059 => sinef <= -8189;
 when 3060 => sinef <= -8190;
 when 3061 => sinef <= -8190;
 when 3062 => sinef <= -8190;
 when 3063 => sinef <= -8190;
 when 3064 => sinef <= -8190;
 when 3065 => sinef <= -8191;
 when 3066 => sinef <= -8191;
 when 3067 => sinef <= -8191;
 when 3068 => sinef <= -8191;
 when 3069 => sinef <= -8191;
 when 3070 => sinef <= -8191;
 when 3071 => sinef <= -8191;
 when 3072 => sinef <= -8191;
 when 3073 => sinef <= -8191;
 when 3074 => sinef <= -8191;
 when 3075 => sinef <= -8191;
 when 3076 => sinef <= -8191;
 when 3077 => sinef <= -8191;
 when 3078 => sinef <= -8191;
 when 3079 => sinef <= -8191;
 when 3080 => sinef <= -8190;
 when 3081 => sinef <= -8190;
 when 3082 => sinef <= -8190;
 when 3083 => sinef <= -8190;
 when 3084 => sinef <= -8190;
 when 3085 => sinef <= -8189;
 when 3086 => sinef <= -8189;
 when 3087 => sinef <= -8189;
 when 3088 => sinef <= -8189;
 when 3089 => sinef <= -8188;
 when 3090 => sinef <= -8188;
 when 3091 => sinef <= -8188;
 when 3092 => sinef <= -8187;
 when 3093 => sinef <= -8187;
 when 3094 => sinef <= -8186;
 when 3095 => sinef <= -8186;
 when 3096 => sinef <= -8185;
 when 3097 => sinef <= -8185;
 when 3098 => sinef <= -8184;
 when 3099 => sinef <= -8184;
 when 3100 => sinef <= -8183;
 when 3101 => sinef <= -8183;
 when 3102 => sinef <= -8182;
 when 3103 => sinef <= -8182;
 when 3104 => sinef <= -8181;
 when 3105 => sinef <= -8181;
 when 3106 => sinef <= -8180;
 when 3107 => sinef <= -8179;
 when 3108 => sinef <= -8179;
 when 3109 => sinef <= -8178;
 when 3110 => sinef <= -8177;
 when 3111 => sinef <= -8176;
 when 3112 => sinef <= -8176;
 when 3113 => sinef <= -8175;
 when 3114 => sinef <= -8174;
 when 3115 => sinef <= -8173;
 when 3116 => sinef <= -8172;
 when 3117 => sinef <= -8171;
 when 3118 => sinef <= -8171;
 when 3119 => sinef <= -8170;
 when 3120 => sinef <= -8169;
 when 3121 => sinef <= -8168;
 when 3122 => sinef <= -8167;
 when 3123 => sinef <= -8166;
 when 3124 => sinef <= -8165;
 when 3125 => sinef <= -8164;
 when 3126 => sinef <= -8163;
 when 3127 => sinef <= -8162;
 when 3128 => sinef <= -8161;
 when 3129 => sinef <= -8160;
 when 3130 => sinef <= -8159;
 when 3131 => sinef <= -8157;
 when 3132 => sinef <= -8156;
 when 3133 => sinef <= -8155;
 when 3134 => sinef <= -8154;
 when 3135 => sinef <= -8153;
 when 3136 => sinef <= -8152;
 when 3137 => sinef <= -8150;
 when 3138 => sinef <= -8149;
 when 3139 => sinef <= -8148;
 when 3140 => sinef <= -8146;
 when 3141 => sinef <= -8145;
 when 3142 => sinef <= -8144;
 when 3143 => sinef <= -8142;
 when 3144 => sinef <= -8141;
 when 3145 => sinef <= -8140;
 when 3146 => sinef <= -8138;
 when 3147 => sinef <= -8137;
 when 3148 => sinef <= -8135;
 when 3149 => sinef <= -8134;
 when 3150 => sinef <= -8132;
 when 3151 => sinef <= -8131;
 when 3152 => sinef <= -8129;
 when 3153 => sinef <= -8128;
 when 3154 => sinef <= -8126;
 when 3155 => sinef <= -8125;
 when 3156 => sinef <= -8123;
 when 3157 => sinef <= -8121;
 when 3158 => sinef <= -8120;
 when 3159 => sinef <= -8118;
 when 3160 => sinef <= -8116;
 when 3161 => sinef <= -8115;
 when 3162 => sinef <= -8113;
 when 3163 => sinef <= -8111;
 when 3164 => sinef <= -8110;
 when 3165 => sinef <= -8108;
 when 3166 => sinef <= -8106;
 when 3167 => sinef <= -8104;
 when 3168 => sinef <= -8102;
 when 3169 => sinef <= -8100;
 when 3170 => sinef <= -8099;
 when 3171 => sinef <= -8097;
 when 3172 => sinef <= -8095;
 when 3173 => sinef <= -8093;
 when 3174 => sinef <= -8091;
 when 3175 => sinef <= -8089;
 when 3176 => sinef <= -8087;
 when 3177 => sinef <= -8085;
 when 3178 => sinef <= -8083;
 when 3179 => sinef <= -8081;
 when 3180 => sinef <= -8079;
 when 3181 => sinef <= -8077;
 when 3182 => sinef <= -8075;
 when 3183 => sinef <= -8073;
 when 3184 => sinef <= -8070;
 when 3185 => sinef <= -8068;
 when 3186 => sinef <= -8066;
 when 3187 => sinef <= -8064;
 when 3188 => sinef <= -8062;
 when 3189 => sinef <= -8059;
 when 3190 => sinef <= -8057;
 when 3191 => sinef <= -8055;
 when 3192 => sinef <= -8053;
 when 3193 => sinef <= -8050;
 when 3194 => sinef <= -8048;
 when 3195 => sinef <= -8046;
 when 3196 => sinef <= -8043;
 when 3197 => sinef <= -8041;
 when 3198 => sinef <= -8038;
 when 3199 => sinef <= -8036;
 when 3200 => sinef <= -8034;
 when 3201 => sinef <= -8031;
 when 3202 => sinef <= -8029;
 when 3203 => sinef <= -8026;
 when 3204 => sinef <= -8024;
 when 3205 => sinef <= -8021;
 when 3206 => sinef <= -8019;
 when 3207 => sinef <= -8016;
 when 3208 => sinef <= -8013;
 when 3209 => sinef <= -8011;
 when 3210 => sinef <= -8008;
 when 3211 => sinef <= -8006;
 when 3212 => sinef <= -8003;
 when 3213 => sinef <= -8000;
 when 3214 => sinef <= -7997;
 when 3215 => sinef <= -7995;
 when 3216 => sinef <= -7992;
 when 3217 => sinef <= -7989;
 when 3218 => sinef <= -7986;
 when 3219 => sinef <= -7984;
 when 3220 => sinef <= -7981;
 when 3221 => sinef <= -7978;
 when 3222 => sinef <= -7975;
 when 3223 => sinef <= -7972;
 when 3224 => sinef <= -7969;
 when 3225 => sinef <= -7966;
 when 3226 => sinef <= -7964;
 when 3227 => sinef <= -7961;
 when 3228 => sinef <= -7958;
 when 3229 => sinef <= -7955;
 when 3230 => sinef <= -7952;
 when 3231 => sinef <= -7949;
 when 3232 => sinef <= -7946;
 when 3233 => sinef <= -7942;
 when 3234 => sinef <= -7939;
 when 3235 => sinef <= -7936;
 when 3236 => sinef <= -7933;
 when 3237 => sinef <= -7930;
 when 3238 => sinef <= -7927;
 when 3239 => sinef <= -7924;
 when 3240 => sinef <= -7921;
 when 3241 => sinef <= -7917;
 when 3242 => sinef <= -7914;
 when 3243 => sinef <= -7911;
 when 3244 => sinef <= -7908;
 when 3245 => sinef <= -7904;
 when 3246 => sinef <= -7901;
 when 3247 => sinef <= -7898;
 when 3248 => sinef <= -7894;
 when 3249 => sinef <= -7891;
 when 3250 => sinef <= -7888;
 when 3251 => sinef <= -7884;
 when 3252 => sinef <= -7881;
 when 3253 => sinef <= -7877;
 when 3254 => sinef <= -7874;
 when 3255 => sinef <= -7870;
 when 3256 => sinef <= -7867;
 when 3257 => sinef <= -7863;
 when 3258 => sinef <= -7860;
 when 3259 => sinef <= -7856;
 when 3260 => sinef <= -7853;
 when 3261 => sinef <= -7849;
 when 3262 => sinef <= -7846;
 when 3263 => sinef <= -7842;
 when 3264 => sinef <= -7838;
 when 3265 => sinef <= -7835;
 when 3266 => sinef <= -7831;
 when 3267 => sinef <= -7827;
 when 3268 => sinef <= -7824;
 when 3269 => sinef <= -7820;
 when 3270 => sinef <= -7816;
 when 3271 => sinef <= -7812;
 when 3272 => sinef <= -7809;
 when 3273 => sinef <= -7805;
 when 3274 => sinef <= -7801;
 when 3275 => sinef <= -7797;
 when 3276 => sinef <= -7793;
 when 3277 => sinef <= -7789;
 when 3278 => sinef <= -7785;
 when 3279 => sinef <= -7782;
 when 3280 => sinef <= -7778;
 when 3281 => sinef <= -7774;
 when 3282 => sinef <= -7770;
 when 3283 => sinef <= -7766;
 when 3284 => sinef <= -7762;
 when 3285 => sinef <= -7758;
 when 3286 => sinef <= -7754;
 when 3287 => sinef <= -7750;
 when 3288 => sinef <= -7745;
 when 3289 => sinef <= -7741;
 when 3290 => sinef <= -7737;
 when 3291 => sinef <= -7733;
 when 3292 => sinef <= -7729;
 when 3293 => sinef <= -7725;
 when 3294 => sinef <= -7721;
 when 3295 => sinef <= -7716;
 when 3296 => sinef <= -7712;
 when 3297 => sinef <= -7708;
 when 3298 => sinef <= -7704;
 when 3299 => sinef <= -7699;
 when 3300 => sinef <= -7695;
 when 3301 => sinef <= -7691;
 when 3302 => sinef <= -7686;
 when 3303 => sinef <= -7682;
 when 3304 => sinef <= -7678;
 when 3305 => sinef <= -7673;
 when 3306 => sinef <= -7669;
 when 3307 => sinef <= -7665;
 when 3308 => sinef <= -7660;
 when 3309 => sinef <= -7656;
 when 3310 => sinef <= -7651;
 when 3311 => sinef <= -7647;
 when 3312 => sinef <= -7642;
 when 3313 => sinef <= -7638;
 when 3314 => sinef <= -7633;
 when 3315 => sinef <= -7628;
 when 3316 => sinef <= -7624;
 when 3317 => sinef <= -7619;
 when 3318 => sinef <= -7615;
 when 3319 => sinef <= -7610;
 when 3320 => sinef <= -7605;
 when 3321 => sinef <= -7601;
 when 3322 => sinef <= -7596;
 when 3323 => sinef <= -7591;
 when 3324 => sinef <= -7587;
 when 3325 => sinef <= -7582;
 when 3326 => sinef <= -7577;
 when 3327 => sinef <= -7572;
 when 3328 => sinef <= -7567;
 when 3329 => sinef <= -7563;
 when 3330 => sinef <= -7558;
 when 3331 => sinef <= -7553;
 when 3332 => sinef <= -7548;
 when 3333 => sinef <= -7543;
 when 3334 => sinef <= -7538;
 when 3335 => sinef <= -7533;
 when 3336 => sinef <= -7528;
 when 3337 => sinef <= -7524;
 when 3338 => sinef <= -7519;
 when 3339 => sinef <= -7514;
 when 3340 => sinef <= -7509;
 when 3341 => sinef <= -7503;
 when 3342 => sinef <= -7498;
 when 3343 => sinef <= -7493;
 when 3344 => sinef <= -7488;
 when 3345 => sinef <= -7483;
 when 3346 => sinef <= -7478;
 when 3347 => sinef <= -7473;
 when 3348 => sinef <= -7468;
 when 3349 => sinef <= -7463;
 when 3350 => sinef <= -7457;
 when 3351 => sinef <= -7452;
 when 3352 => sinef <= -7447;
 when 3353 => sinef <= -7442;
 when 3354 => sinef <= -7436;
 when 3355 => sinef <= -7431;
 when 3356 => sinef <= -7426;
 when 3357 => sinef <= -7421;
 when 3358 => sinef <= -7415;
 when 3359 => sinef <= -7410;
 when 3360 => sinef <= -7405;
 when 3361 => sinef <= -7399;
 when 3362 => sinef <= -7394;
 when 3363 => sinef <= -7388;
 when 3364 => sinef <= -7383;
 when 3365 => sinef <= -7377;
 when 3366 => sinef <= -7372;
 when 3367 => sinef <= -7367;
 when 3368 => sinef <= -7361;
 when 3369 => sinef <= -7356;
 when 3370 => sinef <= -7350;
 when 3371 => sinef <= -7344;
 when 3372 => sinef <= -7339;
 when 3373 => sinef <= -7333;
 when 3374 => sinef <= -7328;
 when 3375 => sinef <= -7322;
 when 3376 => sinef <= -7316;
 when 3377 => sinef <= -7311;
 when 3378 => sinef <= -7305;
 when 3379 => sinef <= -7299;
 when 3380 => sinef <= -7294;
 when 3381 => sinef <= -7288;
 when 3382 => sinef <= -7282;
 when 3383 => sinef <= -7276;
 when 3384 => sinef <= -7271;
 when 3385 => sinef <= -7265;
 when 3386 => sinef <= -7259;
 when 3387 => sinef <= -7253;
 when 3388 => sinef <= -7247;
 when 3389 => sinef <= -7242;
 when 3390 => sinef <= -7236;
 when 3391 => sinef <= -7230;
 when 3392 => sinef <= -7224;
 when 3393 => sinef <= -7218;
 when 3394 => sinef <= -7212;
 when 3395 => sinef <= -7206;
 when 3396 => sinef <= -7200;
 when 3397 => sinef <= -7194;
 when 3398 => sinef <= -7188;
 when 3399 => sinef <= -7182;
 when 3400 => sinef <= -7176;
 when 3401 => sinef <= -7170;
 when 3402 => sinef <= -7164;
 when 3403 => sinef <= -7158;
 when 3404 => sinef <= -7152;
 when 3405 => sinef <= -7145;
 when 3406 => sinef <= -7139;
 when 3407 => sinef <= -7133;
 when 3408 => sinef <= -7127;
 when 3409 => sinef <= -7121;
 when 3410 => sinef <= -7114;
 when 3411 => sinef <= -7108;
 when 3412 => sinef <= -7102;
 when 3413 => sinef <= -7096;
 when 3414 => sinef <= -7089;
 when 3415 => sinef <= -7083;
 when 3416 => sinef <= -7077;
 when 3417 => sinef <= -7070;
 when 3418 => sinef <= -7064;
 when 3419 => sinef <= -7058;
 when 3420 => sinef <= -7051;
 when 3421 => sinef <= -7045;
 when 3422 => sinef <= -7039;
 when 3423 => sinef <= -7032;
 when 3424 => sinef <= -7026;
 when 3425 => sinef <= -7019;
 when 3426 => sinef <= -7013;
 when 3427 => sinef <= -7006;
 when 3428 => sinef <= -7000;
 when 3429 => sinef <= -6993;
 when 3430 => sinef <= -6987;
 when 3431 => sinef <= -6980;
 when 3432 => sinef <= -6973;
 when 3433 => sinef <= -6967;
 when 3434 => sinef <= -6960;
 when 3435 => sinef <= -6954;
 when 3436 => sinef <= -6947;
 when 3437 => sinef <= -6940;
 when 3438 => sinef <= -6934;
 when 3439 => sinef <= -6927;
 when 3440 => sinef <= -6920;
 when 3441 => sinef <= -6913;
 when 3442 => sinef <= -6907;
 when 3443 => sinef <= -6900;
 when 3444 => sinef <= -6893;
 when 3445 => sinef <= -6886;
 when 3446 => sinef <= -6880;
 when 3447 => sinef <= -6873;
 when 3448 => sinef <= -6866;
 when 3449 => sinef <= -6859;
 when 3450 => sinef <= -6852;
 when 3451 => sinef <= -6845;
 when 3452 => sinef <= -6838;
 when 3453 => sinef <= -6831;
 when 3454 => sinef <= -6824;
 when 3455 => sinef <= -6818;
 when 3456 => sinef <= -6811;
 when 3457 => sinef <= -6804;
 when 3458 => sinef <= -6797;
 when 3459 => sinef <= -6790;
 when 3460 => sinef <= -6783;
 when 3461 => sinef <= -6775;
 when 3462 => sinef <= -6768;
 when 3463 => sinef <= -6761;
 when 3464 => sinef <= -6754;
 when 3465 => sinef <= -6747;
 when 3466 => sinef <= -6740;
 when 3467 => sinef <= -6733;
 when 3468 => sinef <= -6726;
 when 3469 => sinef <= -6718;
 when 3470 => sinef <= -6711;
 when 3471 => sinef <= -6704;
 when 3472 => sinef <= -6697;
 when 3473 => sinef <= -6690;
 when 3474 => sinef <= -6682;
 when 3475 => sinef <= -6675;
 when 3476 => sinef <= -6668;
 when 3477 => sinef <= -6660;
 when 3478 => sinef <= -6653;
 when 3479 => sinef <= -6646;
 when 3480 => sinef <= -6638;
 when 3481 => sinef <= -6631;
 when 3482 => sinef <= -6624;
 when 3483 => sinef <= -6616;
 when 3484 => sinef <= -6609;
 when 3485 => sinef <= -6601;
 when 3486 => sinef <= -6594;
 when 3487 => sinef <= -6587;
 when 3488 => sinef <= -6579;
 when 3489 => sinef <= -6572;
 when 3490 => sinef <= -6564;
 when 3491 => sinef <= -6557;
 when 3492 => sinef <= -6549;
 when 3493 => sinef <= -6541;
 when 3494 => sinef <= -6534;
 when 3495 => sinef <= -6526;
 when 3496 => sinef <= -6519;
 when 3497 => sinef <= -6511;
 when 3498 => sinef <= -6503;
 when 3499 => sinef <= -6496;
 when 3500 => sinef <= -6488;
 when 3501 => sinef <= -6480;
 when 3502 => sinef <= -6473;
 when 3503 => sinef <= -6465;
 when 3504 => sinef <= -6457;
 when 3505 => sinef <= -6450;
 when 3506 => sinef <= -6442;
 when 3507 => sinef <= -6434;
 when 3508 => sinef <= -6426;
 when 3509 => sinef <= -6419;
 when 3510 => sinef <= -6411;
 when 3511 => sinef <= -6403;
 when 3512 => sinef <= -6395;
 when 3513 => sinef <= -6387;
 when 3514 => sinef <= -6379;
 when 3515 => sinef <= -6371;
 when 3516 => sinef <= -6363;
 when 3517 => sinef <= -6356;
 when 3518 => sinef <= -6348;
 when 3519 => sinef <= -6340;
 when 3520 => sinef <= -6332;
 when 3521 => sinef <= -6324;
 when 3522 => sinef <= -6316;
 when 3523 => sinef <= -6308;
 when 3524 => sinef <= -6300;
 when 3525 => sinef <= -6292;
 when 3526 => sinef <= -6284;
 when 3527 => sinef <= -6276;
 when 3528 => sinef <= -6267;
 when 3529 => sinef <= -6259;
 when 3530 => sinef <= -6251;
 when 3531 => sinef <= -6243;
 when 3532 => sinef <= -6235;
 when 3533 => sinef <= -6227;
 when 3534 => sinef <= -6219;
 when 3535 => sinef <= -6210;
 when 3536 => sinef <= -6202;
 when 3537 => sinef <= -6194;
 when 3538 => sinef <= -6186;
 when 3539 => sinef <= -6178;
 when 3540 => sinef <= -6169;
 when 3541 => sinef <= -6161;
 when 3542 => sinef <= -6153;
 when 3543 => sinef <= -6144;
 when 3544 => sinef <= -6136;
 when 3545 => sinef <= -6128;
 when 3546 => sinef <= -6120;
 when 3547 => sinef <= -6111;
 when 3548 => sinef <= -6103;
 when 3549 => sinef <= -6094;
 when 3550 => sinef <= -6086;
 when 3551 => sinef <= -6078;
 when 3552 => sinef <= -6069;
 when 3553 => sinef <= -6061;
 when 3554 => sinef <= -6052;
 when 3555 => sinef <= -6044;
 when 3556 => sinef <= -6035;
 when 3557 => sinef <= -6027;
 when 3558 => sinef <= -6018;
 when 3559 => sinef <= -6010;
 when 3560 => sinef <= -6001;
 when 3561 => sinef <= -5993;
 when 3562 => sinef <= -5984;
 when 3563 => sinef <= -5975;
 when 3564 => sinef <= -5967;
 when 3565 => sinef <= -5958;
 when 3566 => sinef <= -5950;
 when 3567 => sinef <= -5941;
 when 3568 => sinef <= -5932;
 when 3569 => sinef <= -5924;
 when 3570 => sinef <= -5915;
 when 3571 => sinef <= -5906;
 when 3572 => sinef <= -5898;
 when 3573 => sinef <= -5889;
 when 3574 => sinef <= -5880;
 when 3575 => sinef <= -5871;
 when 3576 => sinef <= -5863;
 when 3577 => sinef <= -5854;
 when 3578 => sinef <= -5845;
 when 3579 => sinef <= -5836;
 when 3580 => sinef <= -5827;
 when 3581 => sinef <= -5819;
 when 3582 => sinef <= -5810;
 when 3583 => sinef <= -5801;
 when 3584 => sinef <= -5792;
 when 3585 => sinef <= -5783;
 when 3586 => sinef <= -5774;
 when 3587 => sinef <= -5765;
 when 3588 => sinef <= -5756;
 when 3589 => sinef <= -5747;
 when 3590 => sinef <= -5738;
 when 3591 => sinef <= -5729;
 when 3592 => sinef <= -5720;
 when 3593 => sinef <= -5711;
 when 3594 => sinef <= -5702;
 when 3595 => sinef <= -5693;
 when 3596 => sinef <= -5684;
 when 3597 => sinef <= -5675;
 when 3598 => sinef <= -5666;
 when 3599 => sinef <= -5657;
 when 3600 => sinef <= -5648;
 when 3601 => sinef <= -5639;
 when 3602 => sinef <= -5630;
 when 3603 => sinef <= -5621;
 when 3604 => sinef <= -5612;
 when 3605 => sinef <= -5602;
 when 3606 => sinef <= -5593;
 when 3607 => sinef <= -5584;
 when 3608 => sinef <= -5575;
 when 3609 => sinef <= -5566;
 when 3610 => sinef <= -5556;
 when 3611 => sinef <= -5547;
 when 3612 => sinef <= -5538;
 when 3613 => sinef <= -5529;
 when 3614 => sinef <= -5519;
 when 3615 => sinef <= -5510;
 when 3616 => sinef <= -5501;
 when 3617 => sinef <= -5491;
 when 3618 => sinef <= -5482;
 when 3619 => sinef <= -5473;
 when 3620 => sinef <= -5463;
 when 3621 => sinef <= -5454;
 when 3622 => sinef <= -5445;
 when 3623 => sinef <= -5435;
 when 3624 => sinef <= -5426;
 when 3625 => sinef <= -5416;
 when 3626 => sinef <= -5407;
 when 3627 => sinef <= -5398;
 when 3628 => sinef <= -5388;
 when 3629 => sinef <= -5379;
 when 3630 => sinef <= -5369;
 when 3631 => sinef <= -5360;
 when 3632 => sinef <= -5350;
 when 3633 => sinef <= -5341;
 when 3634 => sinef <= -5331;
 when 3635 => sinef <= -5322;
 when 3636 => sinef <= -5312;
 when 3637 => sinef <= -5302;
 when 3638 => sinef <= -5293;
 when 3639 => sinef <= -5283;
 when 3640 => sinef <= -5274;
 when 3641 => sinef <= -5264;
 when 3642 => sinef <= -5254;
 when 3643 => sinef <= -5245;
 when 3644 => sinef <= -5235;
 when 3645 => sinef <= -5225;
 when 3646 => sinef <= -5216;
 when 3647 => sinef <= -5206;
 when 3648 => sinef <= -5196;
 when 3649 => sinef <= -5187;
 when 3650 => sinef <= -5177;
 when 3651 => sinef <= -5167;
 when 3652 => sinef <= -5157;
 when 3653 => sinef <= -5148;
 when 3654 => sinef <= -5138;
 when 3655 => sinef <= -5128;
 when 3656 => sinef <= -5118;
 when 3657 => sinef <= -5108;
 when 3658 => sinef <= -5099;
 when 3659 => sinef <= -5089;
 when 3660 => sinef <= -5079;
 when 3661 => sinef <= -5069;
 when 3662 => sinef <= -5059;
 when 3663 => sinef <= -5049;
 when 3664 => sinef <= -5039;
 when 3665 => sinef <= -5029;
 when 3666 => sinef <= -5020;
 when 3667 => sinef <= -5010;
 when 3668 => sinef <= -5000;
 when 3669 => sinef <= -4990;
 when 3670 => sinef <= -4980;
 when 3671 => sinef <= -4970;
 when 3672 => sinef <= -4960;
 when 3673 => sinef <= -4950;
 when 3674 => sinef <= -4940;
 when 3675 => sinef <= -4930;
 when 3676 => sinef <= -4920;
 when 3677 => sinef <= -4910;
 when 3678 => sinef <= -4900;
 when 3679 => sinef <= -4889;
 when 3680 => sinef <= -4879;
 when 3681 => sinef <= -4869;
 when 3682 => sinef <= -4859;
 when 3683 => sinef <= -4849;
 when 3684 => sinef <= -4839;
 when 3685 => sinef <= -4829;
 when 3686 => sinef <= -4819;
 when 3687 => sinef <= -4808;
 when 3688 => sinef <= -4798;
 when 3689 => sinef <= -4788;
 when 3690 => sinef <= -4778;
 when 3691 => sinef <= -4768;
 when 3692 => sinef <= -4757;
 when 3693 => sinef <= -4747;
 when 3694 => sinef <= -4737;
 when 3695 => sinef <= -4727;
 when 3696 => sinef <= -4716;
 when 3697 => sinef <= -4706;
 when 3698 => sinef <= -4696;
 when 3699 => sinef <= -4686;
 when 3700 => sinef <= -4675;
 when 3701 => sinef <= -4665;
 when 3702 => sinef <= -4655;
 when 3703 => sinef <= -4644;
 when 3704 => sinef <= -4634;
 when 3705 => sinef <= -4624;
 when 3706 => sinef <= -4613;
 when 3707 => sinef <= -4603;
 when 3708 => sinef <= -4592;
 when 3709 => sinef <= -4582;
 when 3710 => sinef <= -4572;
 when 3711 => sinef <= -4561;
 when 3712 => sinef <= -4551;
 when 3713 => sinef <= -4540;
 when 3714 => sinef <= -4530;
 when 3715 => sinef <= -4519;
 when 3716 => sinef <= -4509;
 when 3717 => sinef <= -4498;
 when 3718 => sinef <= -4488;
 when 3719 => sinef <= -4477;
 when 3720 => sinef <= -4467;
 when 3721 => sinef <= -4456;
 when 3722 => sinef <= -4446;
 when 3723 => sinef <= -4435;
 when 3724 => sinef <= -4425;
 when 3725 => sinef <= -4414;
 when 3726 => sinef <= -4403;
 when 3727 => sinef <= -4393;
 when 3728 => sinef <= -4382;
 when 3729 => sinef <= -4372;
 when 3730 => sinef <= -4361;
 when 3731 => sinef <= -4350;
 when 3732 => sinef <= -4340;
 when 3733 => sinef <= -4329;
 when 3734 => sinef <= -4318;
 when 3735 => sinef <= -4308;
 when 3736 => sinef <= -4297;
 when 3737 => sinef <= -4286;
 when 3738 => sinef <= -4275;
 when 3739 => sinef <= -4265;
 when 3740 => sinef <= -4254;
 when 3741 => sinef <= -4243;
 when 3742 => sinef <= -4233;
 when 3743 => sinef <= -4222;
 when 3744 => sinef <= -4211;
 when 3745 => sinef <= -4200;
 when 3746 => sinef <= -4189;
 when 3747 => sinef <= -4179;
 when 3748 => sinef <= -4168;
 when 3749 => sinef <= -4157;
 when 3750 => sinef <= -4146;
 when 3751 => sinef <= -4135;
 when 3752 => sinef <= -4124;
 when 3753 => sinef <= -4114;
 when 3754 => sinef <= -4103;
 when 3755 => sinef <= -4092;
 when 3756 => sinef <= -4081;
 when 3757 => sinef <= -4070;
 when 3758 => sinef <= -4059;
 when 3759 => sinef <= -4048;
 when 3760 => sinef <= -4037;
 when 3761 => sinef <= -4026;
 when 3762 => sinef <= -4015;
 when 3763 => sinef <= -4004;
 when 3764 => sinef <= -3994;
 when 3765 => sinef <= -3983;
 when 3766 => sinef <= -3972;
 when 3767 => sinef <= -3961;
 when 3768 => sinef <= -3950;
 when 3769 => sinef <= -3939;
 when 3770 => sinef <= -3928;
 when 3771 => sinef <= -3917;
 when 3772 => sinef <= -3905;
 when 3773 => sinef <= -3894;
 when 3774 => sinef <= -3883;
 when 3775 => sinef <= -3872;
 when 3776 => sinef <= -3861;
 when 3777 => sinef <= -3850;
 when 3778 => sinef <= -3839;
 when 3779 => sinef <= -3828;
 when 3780 => sinef <= -3817;
 when 3781 => sinef <= -3806;
 when 3782 => sinef <= -3795;
 when 3783 => sinef <= -3783;
 when 3784 => sinef <= -3772;
 when 3785 => sinef <= -3761;
 when 3786 => sinef <= -3750;
 when 3787 => sinef <= -3739;
 when 3788 => sinef <= -3728;
 when 3789 => sinef <= -3716;
 when 3790 => sinef <= -3705;
 when 3791 => sinef <= -3694;
 when 3792 => sinef <= -3683;
 when 3793 => sinef <= -3672;
 when 3794 => sinef <= -3660;
 when 3795 => sinef <= -3649;
 when 3796 => sinef <= -3638;
 when 3797 => sinef <= -3627;
 when 3798 => sinef <= -3615;
 when 3799 => sinef <= -3604;
 when 3800 => sinef <= -3593;
 when 3801 => sinef <= -3581;
 when 3802 => sinef <= -3570;
 when 3803 => sinef <= -3559;
 when 3804 => sinef <= -3547;
 when 3805 => sinef <= -3536;
 when 3806 => sinef <= -3525;
 when 3807 => sinef <= -3513;
 when 3808 => sinef <= -3502;
 when 3809 => sinef <= -3491;
 when 3810 => sinef <= -3479;
 when 3811 => sinef <= -3468;
 when 3812 => sinef <= -3457;
 when 3813 => sinef <= -3445;
 when 3814 => sinef <= -3434;
 when 3815 => sinef <= -3422;
 when 3816 => sinef <= -3411;
 when 3817 => sinef <= -3400;
 when 3818 => sinef <= -3388;
 when 3819 => sinef <= -3377;
 when 3820 => sinef <= -3365;
 when 3821 => sinef <= -3354;
 when 3822 => sinef <= -3342;
 when 3823 => sinef <= -3331;
 when 3824 => sinef <= -3319;
 when 3825 => sinef <= -3308;
 when 3826 => sinef <= -3296;
 when 3827 => sinef <= -3285;
 when 3828 => sinef <= -3273;
 when 3829 => sinef <= -3262;
 when 3830 => sinef <= -3250;
 when 3831 => sinef <= -3239;
 when 3832 => sinef <= -3227;
 when 3833 => sinef <= -3216;
 when 3834 => sinef <= -3204;
 when 3835 => sinef <= -3193;
 when 3836 => sinef <= -3181;
 when 3837 => sinef <= -3169;
 when 3838 => sinef <= -3158;
 when 3839 => sinef <= -3146;
 when 3840 => sinef <= -3135;
 when 3841 => sinef <= -3123;
 when 3842 => sinef <= -3111;
 when 3843 => sinef <= -3100;
 when 3844 => sinef <= -3088;
 when 3845 => sinef <= -3076;
 when 3846 => sinef <= -3065;
 when 3847 => sinef <= -3053;
 when 3848 => sinef <= -3041;
 when 3849 => sinef <= -3030;
 when 3850 => sinef <= -3018;
 when 3851 => sinef <= -3006;
 when 3852 => sinef <= -2995;
 when 3853 => sinef <= -2983;
 when 3854 => sinef <= -2971;
 when 3855 => sinef <= -2960;
 when 3856 => sinef <= -2948;
 when 3857 => sinef <= -2936;
 when 3858 => sinef <= -2924;
 when 3859 => sinef <= -2913;
 when 3860 => sinef <= -2901;
 when 3861 => sinef <= -2889;
 when 3862 => sinef <= -2877;
 when 3863 => sinef <= -2866;
 when 3864 => sinef <= -2854;
 when 3865 => sinef <= -2842;
 when 3866 => sinef <= -2830;
 when 3867 => sinef <= -2819;
 when 3868 => sinef <= -2807;
 when 3869 => sinef <= -2795;
 when 3870 => sinef <= -2783;
 when 3871 => sinef <= -2771;
 when 3872 => sinef <= -2759;
 when 3873 => sinef <= -2748;
 when 3874 => sinef <= -2736;
 when 3875 => sinef <= -2724;
 when 3876 => sinef <= -2712;
 when 3877 => sinef <= -2700;
 when 3878 => sinef <= -2688;
 when 3879 => sinef <= -2676;
 when 3880 => sinef <= -2665;
 when 3881 => sinef <= -2653;
 when 3882 => sinef <= -2641;
 when 3883 => sinef <= -2629;
 when 3884 => sinef <= -2617;
 when 3885 => sinef <= -2605;
 when 3886 => sinef <= -2593;
 when 3887 => sinef <= -2581;
 when 3888 => sinef <= -2569;
 when 3889 => sinef <= -2557;
 when 3890 => sinef <= -2545;
 when 3891 => sinef <= -2534;
 when 3892 => sinef <= -2522;
 when 3893 => sinef <= -2510;
 when 3894 => sinef <= -2498;
 when 3895 => sinef <= -2486;
 when 3896 => sinef <= -2474;
 when 3897 => sinef <= -2462;
 when 3898 => sinef <= -2450;
 when 3899 => sinef <= -2438;
 when 3900 => sinef <= -2426;
 when 3901 => sinef <= -2414;
 when 3902 => sinef <= -2402;
 when 3903 => sinef <= -2390;
 when 3904 => sinef <= -2378;
 when 3905 => sinef <= -2366;
 when 3906 => sinef <= -2354;
 when 3907 => sinef <= -2342;
 when 3908 => sinef <= -2330;
 when 3909 => sinef <= -2318;
 when 3910 => sinef <= -2305;
 when 3911 => sinef <= -2293;
 when 3912 => sinef <= -2281;
 when 3913 => sinef <= -2269;
 when 3914 => sinef <= -2257;
 when 3915 => sinef <= -2245;
 when 3916 => sinef <= -2233;
 when 3917 => sinef <= -2221;
 when 3918 => sinef <= -2209;
 when 3919 => sinef <= -2197;
 when 3920 => sinef <= -2185;
 when 3921 => sinef <= -2173;
 when 3922 => sinef <= -2160;
 when 3923 => sinef <= -2148;
 when 3924 => sinef <= -2136;
 when 3925 => sinef <= -2124;
 when 3926 => sinef <= -2112;
 when 3927 => sinef <= -2100;
 when 3928 => sinef <= -2088;
 when 3929 => sinef <= -2075;
 when 3930 => sinef <= -2063;
 when 3931 => sinef <= -2051;
 when 3932 => sinef <= -2039;
 when 3933 => sinef <= -2027;
 when 3934 => sinef <= -2015;
 when 3935 => sinef <= -2002;
 when 3936 => sinef <= -1990;
 when 3937 => sinef <= -1978;
 when 3938 => sinef <= -1966;
 when 3939 => sinef <= -1954;
 when 3940 => sinef <= -1941;
 when 3941 => sinef <= -1929;
 when 3942 => sinef <= -1917;
 when 3943 => sinef <= -1905;
 when 3944 => sinef <= -1893;
 when 3945 => sinef <= -1880;
 when 3946 => sinef <= -1868;
 when 3947 => sinef <= -1856;
 when 3948 => sinef <= -1844;
 when 3949 => sinef <= -1831;
 when 3950 => sinef <= -1819;
 when 3951 => sinef <= -1807;
 when 3952 => sinef <= -1795;
 when 3953 => sinef <= -1782;
 when 3954 => sinef <= -1770;
 when 3955 => sinef <= -1758;
 when 3956 => sinef <= -1746;
 when 3957 => sinef <= -1733;
 when 3958 => sinef <= -1721;
 when 3959 => sinef <= -1709;
 when 3960 => sinef <= -1696;
 when 3961 => sinef <= -1684;
 when 3962 => sinef <= -1672;
 when 3963 => sinef <= -1660;
 when 3964 => sinef <= -1647;
 when 3965 => sinef <= -1635;
 when 3966 => sinef <= -1623;
 when 3967 => sinef <= -1610;
 when 3968 => sinef <= -1598;
 when 3969 => sinef <= -1586;
 when 3970 => sinef <= -1573;
 when 3971 => sinef <= -1561;
 when 3972 => sinef <= -1549;
 when 3973 => sinef <= -1536;
 when 3974 => sinef <= -1524;
 when 3975 => sinef <= -1512;
 when 3976 => sinef <= -1499;
 when 3977 => sinef <= -1487;
 when 3978 => sinef <= -1475;
 when 3979 => sinef <= -1462;
 when 3980 => sinef <= -1450;
 when 3981 => sinef <= -1437;
 when 3982 => sinef <= -1425;
 when 3983 => sinef <= -1413;
 when 3984 => sinef <= -1400;
 when 3985 => sinef <= -1388;
 when 3986 => sinef <= -1376;
 when 3987 => sinef <= -1363;
 when 3988 => sinef <= -1351;
 when 3989 => sinef <= -1338;
 when 3990 => sinef <= -1326;
 when 3991 => sinef <= -1314;
 when 3992 => sinef <= -1301;
 when 3993 => sinef <= -1289;
 when 3994 => sinef <= -1276;
 when 3995 => sinef <= -1264;
 when 3996 => sinef <= -1252;
 when 3997 => sinef <= -1239;
 when 3998 => sinef <= -1227;
 when 3999 => sinef <= -1214;
 when 4000 => sinef <= -1202;
 when 4001 => sinef <= -1189;
 when 4002 => sinef <= -1177;
 when 4003 => sinef <= -1165;
 when 4004 => sinef <= -1152;
 when 4005 => sinef <= -1140;
 when 4006 => sinef <= -1127;
 when 4007 => sinef <= -1115;
 when 4008 => sinef <= -1102;
 when 4009 => sinef <= -1090;
 when 4010 => sinef <= -1077;
 when 4011 => sinef <= -1065;
 when 4012 => sinef <= -1053;
 when 4013 => sinef <= -1040;
 when 4014 => sinef <= -1028;
 when 4015 => sinef <= -1015;
 when 4016 => sinef <= -1003;
 when 4017 => sinef <= -990;
 when 4018 => sinef <= -978;
 when 4019 => sinef <= -965;
 when 4020 => sinef <= -953;
 when 4021 => sinef <= -940;
 when 4022 => sinef <= -928;
 when 4023 => sinef <= -915;
 when 4024 => sinef <= -903;
 when 4025 => sinef <= -890;
 when 4026 => sinef <= -878;
 when 4027 => sinef <= -865;
 when 4028 => sinef <= -853;
 when 4029 => sinef <= -840;
 when 4030 => sinef <= -828;
 when 4031 => sinef <= -815;
 when 4032 => sinef <= -803;
 when 4033 => sinef <= -790;
 when 4034 => sinef <= -778;
 when 4035 => sinef <= -765;
 when 4036 => sinef <= -753;
 when 4037 => sinef <= -740;
 when 4038 => sinef <= -728;
 when 4039 => sinef <= -715;
 when 4040 => sinef <= -703;
 when 4041 => sinef <= -690;
 when 4042 => sinef <= -678;
 when 4043 => sinef <= -665;
 when 4044 => sinef <= -653;
 when 4045 => sinef <= -640;
 when 4046 => sinef <= -628;
 when 4047 => sinef <= -615;
 when 4048 => sinef <= -603;
 when 4049 => sinef <= -590;
 when 4050 => sinef <= -578;
 when 4051 => sinef <= -565;
 when 4052 => sinef <= -552;
 when 4053 => sinef <= -540;
 when 4054 => sinef <= -527;
 when 4055 => sinef <= -515;
 when 4056 => sinef <= -502;
 when 4057 => sinef <= -490;
 when 4058 => sinef <= -477;
 when 4059 => sinef <= -465;
 when 4060 => sinef <= -452;
 when 4061 => sinef <= -440;
 when 4062 => sinef <= -427;
 when 4063 => sinef <= -414;
 when 4064 => sinef <= -402;
 when 4065 => sinef <= -389;
 when 4066 => sinef <= -377;
 when 4067 => sinef <= -364;
 when 4068 => sinef <= -352;
 when 4069 => sinef <= -339;
 when 4070 => sinef <= -327;
 when 4071 => sinef <= -314;
 when 4072 => sinef <= -301;
 when 4073 => sinef <= -289;
 when 4074 => sinef <= -276;
 when 4075 => sinef <= -264;
 when 4076 => sinef <= -251;
 when 4077 => sinef <= -239;
 when 4078 => sinef <= -226;
 when 4079 => sinef <= -214;
 when 4080 => sinef <= -201;
 when 4081 => sinef <= -188;
 when 4082 => sinef <= -176;
 when 4083 => sinef <= -163;
 when 4084 => sinef <= -151;
 when 4085 => sinef <= -138;
 when 4086 => sinef <= -126;
 when 4087 => sinef <= -113;
 when 4088 => sinef <= -101;
 when 4089 => sinef <= -88;
 when 4090 => sinef <= -75;
 when 4091 => sinef <= -63;
 when 4092 => sinef <= -50;
 when 4093 => sinef <= -38;
 when 4094 => sinef <= -25;
 when 4095 => sinef <= -13;
	 when others => sinef <=0;
	end case;
	end if;
end process;
	
	
end rtl;


